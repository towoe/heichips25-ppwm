module heichips25_ppwm (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire \u_ppwm/global_counter[0] ;
 wire \u_ppwm/global_counter[10] ;
 wire \u_ppwm/global_counter[11] ;
 wire \u_ppwm/global_counter[12] ;
 wire \u_ppwm/global_counter[13] ;
 wire \u_ppwm/global_counter[14] ;
 wire \u_ppwm/global_counter[15] ;
 wire \u_ppwm/global_counter[16] ;
 wire \u_ppwm/global_counter[17] ;
 wire \u_ppwm/global_counter[18] ;
 wire \u_ppwm/global_counter[19] ;
 wire \u_ppwm/global_counter[1] ;
 wire \u_ppwm/global_counter[2] ;
 wire \u_ppwm/global_counter[3] ;
 wire \u_ppwm/global_counter[4] ;
 wire \u_ppwm/global_counter[5] ;
 wire \u_ppwm/global_counter[6] ;
 wire \u_ppwm/global_counter[7] ;
 wire \u_ppwm/global_counter[8] ;
 wire \u_ppwm/global_counter[9] ;
 wire \u_ppwm/instr[0] ;
 wire \u_ppwm/instr[1] ;
 wire \u_ppwm/instr[2] ;
 wire \u_ppwm/instr[3] ;
 wire \u_ppwm/instr[4] ;
 wire \u_ppwm/instr[5] ;
 wire \u_ppwm/instr[6] ;
 wire \u_ppwm/mem_write_done ;
 wire \u_ppwm/pc[0] ;
 wire \u_ppwm/pc[1] ;
 wire \u_ppwm/pc[2] ;
 wire \u_ppwm/pc[3] ;
 wire \u_ppwm/period_start ;
 wire \u_ppwm/polarity ;
 wire \u_ppwm/pwm_value[0] ;
 wire \u_ppwm/pwm_value[1] ;
 wire \u_ppwm/pwm_value[2] ;
 wire \u_ppwm/pwm_value[3] ;
 wire \u_ppwm/pwm_value[4] ;
 wire \u_ppwm/pwm_value[5] ;
 wire \u_ppwm/pwm_value[6] ;
 wire \u_ppwm/pwm_value[7] ;
 wire \u_ppwm/pwm_value[8] ;
 wire \u_ppwm/pwm_value[9] ;
 wire \u_ppwm/u_ex/_0000_ ;
 wire \u_ppwm/u_ex/_0001_ ;
 wire \u_ppwm/u_ex/_0002_ ;
 wire \u_ppwm/u_ex/_0003_ ;
 wire \u_ppwm/u_ex/_0004_ ;
 wire \u_ppwm/u_ex/_0005_ ;
 wire \u_ppwm/u_ex/_0006_ ;
 wire \u_ppwm/u_ex/_0007_ ;
 wire \u_ppwm/u_ex/_0008_ ;
 wire \u_ppwm/u_ex/_0009_ ;
 wire \u_ppwm/u_ex/_0010_ ;
 wire \u_ppwm/u_ex/_0011_ ;
 wire \u_ppwm/u_ex/_0012_ ;
 wire \u_ppwm/u_ex/_0013_ ;
 wire \u_ppwm/u_ex/_0014_ ;
 wire \u_ppwm/u_ex/_0015_ ;
 wire \u_ppwm/u_ex/_0016_ ;
 wire \u_ppwm/u_ex/_0017_ ;
 wire \u_ppwm/u_ex/_0018_ ;
 wire \u_ppwm/u_ex/_0019_ ;
 wire \u_ppwm/u_ex/_0020_ ;
 wire \u_ppwm/u_ex/_0021_ ;
 wire \u_ppwm/u_ex/_0022_ ;
 wire \u_ppwm/u_ex/_0023_ ;
 wire \u_ppwm/u_ex/_0024_ ;
 wire \u_ppwm/u_ex/_0025_ ;
 wire \u_ppwm/u_ex/_0026_ ;
 wire \u_ppwm/u_ex/_0027_ ;
 wire \u_ppwm/u_ex/_0028_ ;
 wire \u_ppwm/u_ex/_0029_ ;
 wire \u_ppwm/u_ex/_0030_ ;
 wire \u_ppwm/u_ex/_0031_ ;
 wire \u_ppwm/u_ex/_0032_ ;
 wire \u_ppwm/u_ex/_0033_ ;
 wire \u_ppwm/u_ex/_0034_ ;
 wire \u_ppwm/u_ex/_0035_ ;
 wire \u_ppwm/u_ex/_0036_ ;
 wire \u_ppwm/u_ex/_0037_ ;
 wire \u_ppwm/u_ex/_0038_ ;
 wire \u_ppwm/u_ex/_0039_ ;
 wire \u_ppwm/u_ex/_0040_ ;
 wire \u_ppwm/u_ex/_0041_ ;
 wire \u_ppwm/u_ex/_0042_ ;
 wire \u_ppwm/u_ex/_0043_ ;
 wire \u_ppwm/u_ex/_0044_ ;
 wire \u_ppwm/u_ex/_0045_ ;
 wire \u_ppwm/u_ex/_0046_ ;
 wire \u_ppwm/u_ex/_0047_ ;
 wire \u_ppwm/u_ex/_0048_ ;
 wire \u_ppwm/u_ex/_0049_ ;
 wire \u_ppwm/u_ex/_0050_ ;
 wire \u_ppwm/u_ex/_0051_ ;
 wire \u_ppwm/u_ex/_0052_ ;
 wire \u_ppwm/u_ex/_0053_ ;
 wire \u_ppwm/u_ex/_0054_ ;
 wire \u_ppwm/u_ex/_0055_ ;
 wire \u_ppwm/u_ex/_0056_ ;
 wire \u_ppwm/u_ex/_0057_ ;
 wire \u_ppwm/u_ex/_0058_ ;
 wire \u_ppwm/u_ex/_0059_ ;
 wire \u_ppwm/u_ex/_0060_ ;
 wire \u_ppwm/u_ex/_0061_ ;
 wire \u_ppwm/u_ex/_0062_ ;
 wire \u_ppwm/u_ex/_0063_ ;
 wire \u_ppwm/u_ex/_0064_ ;
 wire \u_ppwm/u_ex/_0065_ ;
 wire \u_ppwm/u_ex/_0066_ ;
 wire \u_ppwm/u_ex/_0067_ ;
 wire \u_ppwm/u_ex/_0068_ ;
 wire \u_ppwm/u_ex/_0069_ ;
 wire \u_ppwm/u_ex/_0070_ ;
 wire \u_ppwm/u_ex/_0071_ ;
 wire \u_ppwm/u_ex/_0072_ ;
 wire \u_ppwm/u_ex/_0073_ ;
 wire \u_ppwm/u_ex/_0074_ ;
 wire \u_ppwm/u_ex/_0075_ ;
 wire \u_ppwm/u_ex/_0076_ ;
 wire \u_ppwm/u_ex/_0077_ ;
 wire \u_ppwm/u_ex/_0078_ ;
 wire \u_ppwm/u_ex/_0079_ ;
 wire \u_ppwm/u_ex/_0080_ ;
 wire \u_ppwm/u_ex/_0081_ ;
 wire \u_ppwm/u_ex/_0082_ ;
 wire \u_ppwm/u_ex/_0083_ ;
 wire \u_ppwm/u_ex/_0084_ ;
 wire \u_ppwm/u_ex/_0085_ ;
 wire \u_ppwm/u_ex/_0086_ ;
 wire \u_ppwm/u_ex/_0087_ ;
 wire \u_ppwm/u_ex/_0088_ ;
 wire \u_ppwm/u_ex/_0089_ ;
 wire \u_ppwm/u_ex/_0090_ ;
 wire \u_ppwm/u_ex/_0091_ ;
 wire \u_ppwm/u_ex/_0092_ ;
 wire \u_ppwm/u_ex/_0093_ ;
 wire \u_ppwm/u_ex/_0094_ ;
 wire \u_ppwm/u_ex/_0095_ ;
 wire \u_ppwm/u_ex/_0096_ ;
 wire \u_ppwm/u_ex/_0097_ ;
 wire \u_ppwm/u_ex/_0098_ ;
 wire \u_ppwm/u_ex/_0099_ ;
 wire \u_ppwm/u_ex/_0100_ ;
 wire \u_ppwm/u_ex/_0101_ ;
 wire \u_ppwm/u_ex/_0102_ ;
 wire \u_ppwm/u_ex/_0103_ ;
 wire \u_ppwm/u_ex/_0104_ ;
 wire \u_ppwm/u_ex/_0105_ ;
 wire \u_ppwm/u_ex/_0106_ ;
 wire \u_ppwm/u_ex/_0107_ ;
 wire \u_ppwm/u_ex/_0108_ ;
 wire \u_ppwm/u_ex/_0109_ ;
 wire \u_ppwm/u_ex/_0110_ ;
 wire \u_ppwm/u_ex/_0111_ ;
 wire \u_ppwm/u_ex/_0112_ ;
 wire \u_ppwm/u_ex/_0113_ ;
 wire \u_ppwm/u_ex/_0114_ ;
 wire \u_ppwm/u_ex/_0115_ ;
 wire \u_ppwm/u_ex/_0116_ ;
 wire \u_ppwm/u_ex/_0117_ ;
 wire \u_ppwm/u_ex/_0118_ ;
 wire \u_ppwm/u_ex/_0119_ ;
 wire \u_ppwm/u_ex/_0120_ ;
 wire \u_ppwm/u_ex/_0121_ ;
 wire \u_ppwm/u_ex/_0122_ ;
 wire \u_ppwm/u_ex/_0123_ ;
 wire \u_ppwm/u_ex/_0124_ ;
 wire \u_ppwm/u_ex/_0125_ ;
 wire \u_ppwm/u_ex/_0126_ ;
 wire \u_ppwm/u_ex/_0127_ ;
 wire \u_ppwm/u_ex/_0128_ ;
 wire \u_ppwm/u_ex/_0129_ ;
 wire \u_ppwm/u_ex/_0130_ ;
 wire \u_ppwm/u_ex/_0131_ ;
 wire \u_ppwm/u_ex/_0132_ ;
 wire \u_ppwm/u_ex/_0133_ ;
 wire \u_ppwm/u_ex/_0134_ ;
 wire \u_ppwm/u_ex/_0135_ ;
 wire \u_ppwm/u_ex/_0136_ ;
 wire \u_ppwm/u_ex/_0137_ ;
 wire \u_ppwm/u_ex/_0138_ ;
 wire \u_ppwm/u_ex/_0139_ ;
 wire \u_ppwm/u_ex/_0140_ ;
 wire \u_ppwm/u_ex/_0141_ ;
 wire \u_ppwm/u_ex/_0142_ ;
 wire \u_ppwm/u_ex/_0143_ ;
 wire \u_ppwm/u_ex/_0144_ ;
 wire \u_ppwm/u_ex/_0145_ ;
 wire \u_ppwm/u_ex/_0146_ ;
 wire \u_ppwm/u_ex/_0147_ ;
 wire \u_ppwm/u_ex/_0148_ ;
 wire \u_ppwm/u_ex/_0149_ ;
 wire \u_ppwm/u_ex/_0150_ ;
 wire \u_ppwm/u_ex/_0151_ ;
 wire \u_ppwm/u_ex/_0152_ ;
 wire \u_ppwm/u_ex/_0153_ ;
 wire \u_ppwm/u_ex/_0154_ ;
 wire \u_ppwm/u_ex/_0155_ ;
 wire \u_ppwm/u_ex/_0156_ ;
 wire \u_ppwm/u_ex/_0157_ ;
 wire \u_ppwm/u_ex/_0158_ ;
 wire \u_ppwm/u_ex/_0159_ ;
 wire \u_ppwm/u_ex/_0160_ ;
 wire \u_ppwm/u_ex/_0161_ ;
 wire \u_ppwm/u_ex/_0162_ ;
 wire \u_ppwm/u_ex/_0163_ ;
 wire \u_ppwm/u_ex/_0164_ ;
 wire \u_ppwm/u_ex/_0165_ ;
 wire \u_ppwm/u_ex/_0166_ ;
 wire \u_ppwm/u_ex/_0167_ ;
 wire \u_ppwm/u_ex/_0168_ ;
 wire \u_ppwm/u_ex/_0169_ ;
 wire \u_ppwm/u_ex/_0170_ ;
 wire \u_ppwm/u_ex/_0171_ ;
 wire \u_ppwm/u_ex/_0172_ ;
 wire \u_ppwm/u_ex/_0173_ ;
 wire \u_ppwm/u_ex/_0174_ ;
 wire \u_ppwm/u_ex/_0175_ ;
 wire \u_ppwm/u_ex/_0176_ ;
 wire \u_ppwm/u_ex/_0177_ ;
 wire \u_ppwm/u_ex/_0178_ ;
 wire \u_ppwm/u_ex/_0179_ ;
 wire \u_ppwm/u_ex/_0180_ ;
 wire \u_ppwm/u_ex/_0181_ ;
 wire \u_ppwm/u_ex/_0182_ ;
 wire \u_ppwm/u_ex/_0183_ ;
 wire \u_ppwm/u_ex/_0184_ ;
 wire \u_ppwm/u_ex/_0185_ ;
 wire \u_ppwm/u_ex/_0186_ ;
 wire \u_ppwm/u_ex/_0187_ ;
 wire \u_ppwm/u_ex/_0188_ ;
 wire \u_ppwm/u_ex/_0189_ ;
 wire \u_ppwm/u_ex/_0190_ ;
 wire \u_ppwm/u_ex/_0191_ ;
 wire \u_ppwm/u_ex/_0192_ ;
 wire \u_ppwm/u_ex/_0193_ ;
 wire \u_ppwm/u_ex/_0194_ ;
 wire \u_ppwm/u_ex/_0195_ ;
 wire \u_ppwm/u_ex/_0196_ ;
 wire \u_ppwm/u_ex/_0197_ ;
 wire \u_ppwm/u_ex/_0198_ ;
 wire \u_ppwm/u_ex/_0199_ ;
 wire \u_ppwm/u_ex/_0200_ ;
 wire \u_ppwm/u_ex/_0201_ ;
 wire \u_ppwm/u_ex/_0202_ ;
 wire \u_ppwm/u_ex/_0203_ ;
 wire \u_ppwm/u_ex/_0204_ ;
 wire \u_ppwm/u_ex/_0205_ ;
 wire \u_ppwm/u_ex/_0206_ ;
 wire \u_ppwm/u_ex/_0207_ ;
 wire \u_ppwm/u_ex/_0208_ ;
 wire \u_ppwm/u_ex/_0209_ ;
 wire \u_ppwm/u_ex/_0210_ ;
 wire \u_ppwm/u_ex/_0211_ ;
 wire \u_ppwm/u_ex/_0212_ ;
 wire \u_ppwm/u_ex/_0213_ ;
 wire \u_ppwm/u_ex/_0214_ ;
 wire \u_ppwm/u_ex/_0215_ ;
 wire \u_ppwm/u_ex/_0216_ ;
 wire \u_ppwm/u_ex/_0217_ ;
 wire \u_ppwm/u_ex/_0218_ ;
 wire \u_ppwm/u_ex/_0219_ ;
 wire \u_ppwm/u_ex/_0220_ ;
 wire \u_ppwm/u_ex/_0221_ ;
 wire \u_ppwm/u_ex/_0222_ ;
 wire \u_ppwm/u_ex/_0223_ ;
 wire \u_ppwm/u_ex/_0224_ ;
 wire \u_ppwm/u_ex/_0225_ ;
 wire \u_ppwm/u_ex/_0226_ ;
 wire \u_ppwm/u_ex/_0227_ ;
 wire \u_ppwm/u_ex/_0228_ ;
 wire \u_ppwm/u_ex/_0229_ ;
 wire \u_ppwm/u_ex/_0230_ ;
 wire \u_ppwm/u_ex/_0231_ ;
 wire \u_ppwm/u_ex/_0232_ ;
 wire \u_ppwm/u_ex/_0233_ ;
 wire \u_ppwm/u_ex/_0234_ ;
 wire \u_ppwm/u_ex/_0235_ ;
 wire \u_ppwm/u_ex/_0236_ ;
 wire \u_ppwm/u_ex/_0237_ ;
 wire \u_ppwm/u_ex/_0238_ ;
 wire \u_ppwm/u_ex/_0239_ ;
 wire \u_ppwm/u_ex/_0240_ ;
 wire \u_ppwm/u_ex/_0241_ ;
 wire \u_ppwm/u_ex/_0242_ ;
 wire \u_ppwm/u_ex/_0243_ ;
 wire \u_ppwm/u_ex/_0244_ ;
 wire \u_ppwm/u_ex/_0245_ ;
 wire \u_ppwm/u_ex/_0246_ ;
 wire \u_ppwm/u_ex/_0247_ ;
 wire \u_ppwm/u_ex/_0248_ ;
 wire \u_ppwm/u_ex/_0249_ ;
 wire \u_ppwm/u_ex/_0250_ ;
 wire \u_ppwm/u_ex/_0251_ ;
 wire \u_ppwm/u_ex/_0252_ ;
 wire \u_ppwm/u_ex/_0253_ ;
 wire \u_ppwm/u_ex/_0254_ ;
 wire \u_ppwm/u_ex/_0255_ ;
 wire \u_ppwm/u_ex/_0256_ ;
 wire \u_ppwm/u_ex/_0257_ ;
 wire \u_ppwm/u_ex/_0258_ ;
 wire \u_ppwm/u_ex/_0259_ ;
 wire \u_ppwm/u_ex/_0260_ ;
 wire \u_ppwm/u_ex/_0261_ ;
 wire \u_ppwm/u_ex/_0262_ ;
 wire \u_ppwm/u_ex/_0263_ ;
 wire \u_ppwm/u_ex/_0264_ ;
 wire \u_ppwm/u_ex/_0265_ ;
 wire \u_ppwm/u_ex/_0266_ ;
 wire \u_ppwm/u_ex/_0267_ ;
 wire \u_ppwm/u_ex/_0268_ ;
 wire \u_ppwm/u_ex/_0269_ ;
 wire \u_ppwm/u_ex/_0270_ ;
 wire \u_ppwm/u_ex/_0271_ ;
 wire \u_ppwm/u_ex/_0272_ ;
 wire \u_ppwm/u_ex/_0273_ ;
 wire \u_ppwm/u_ex/_0274_ ;
 wire \u_ppwm/u_ex/_0275_ ;
 wire \u_ppwm/u_ex/_0276_ ;
 wire \u_ppwm/u_ex/_0277_ ;
 wire \u_ppwm/u_ex/_0278_ ;
 wire \u_ppwm/u_ex/_0279_ ;
 wire \u_ppwm/u_ex/_0280_ ;
 wire \u_ppwm/u_ex/_0281_ ;
 wire \u_ppwm/u_ex/_0282_ ;
 wire \u_ppwm/u_ex/_0283_ ;
 wire \u_ppwm/u_ex/_0284_ ;
 wire \u_ppwm/u_ex/_0285_ ;
 wire \u_ppwm/u_ex/_0286_ ;
 wire \u_ppwm/u_ex/_0287_ ;
 wire \u_ppwm/u_ex/_0288_ ;
 wire \u_ppwm/u_ex/_0289_ ;
 wire \u_ppwm/u_ex/_0290_ ;
 wire \u_ppwm/u_ex/_0291_ ;
 wire \u_ppwm/u_ex/_0292_ ;
 wire \u_ppwm/u_ex/_0293_ ;
 wire \u_ppwm/u_ex/_0294_ ;
 wire \u_ppwm/u_ex/_0295_ ;
 wire \u_ppwm/u_ex/_0296_ ;
 wire \u_ppwm/u_ex/_0297_ ;
 wire \u_ppwm/u_ex/_0298_ ;
 wire \u_ppwm/u_ex/_0299_ ;
 wire \u_ppwm/u_ex/_0300_ ;
 wire \u_ppwm/u_ex/_0301_ ;
 wire \u_ppwm/u_ex/_0302_ ;
 wire \u_ppwm/u_ex/_0303_ ;
 wire \u_ppwm/u_ex/_0304_ ;
 wire \u_ppwm/u_ex/_0305_ ;
 wire \u_ppwm/u_ex/_0306_ ;
 wire \u_ppwm/u_ex/_0307_ ;
 wire \u_ppwm/u_ex/_0308_ ;
 wire \u_ppwm/u_ex/_0309_ ;
 wire \u_ppwm/u_ex/_0310_ ;
 wire \u_ppwm/u_ex/_0311_ ;
 wire \u_ppwm/u_ex/_0312_ ;
 wire \u_ppwm/u_ex/_0313_ ;
 wire \u_ppwm/u_ex/_0314_ ;
 wire \u_ppwm/u_ex/_0315_ ;
 wire \u_ppwm/u_ex/_0316_ ;
 wire \u_ppwm/u_ex/_0317_ ;
 wire \u_ppwm/u_ex/_0318_ ;
 wire \u_ppwm/u_ex/_0319_ ;
 wire \u_ppwm/u_ex/_0320_ ;
 wire \u_ppwm/u_ex/_0321_ ;
 wire \u_ppwm/u_ex/_0322_ ;
 wire \u_ppwm/u_ex/_0323_ ;
 wire \u_ppwm/u_ex/_0324_ ;
 wire \u_ppwm/u_ex/_0325_ ;
 wire \u_ppwm/u_ex/_0326_ ;
 wire \u_ppwm/u_ex/_0327_ ;
 wire \u_ppwm/u_ex/_0328_ ;
 wire \u_ppwm/u_ex/_0329_ ;
 wire \u_ppwm/u_ex/_0330_ ;
 wire \u_ppwm/u_ex/_0331_ ;
 wire \u_ppwm/u_ex/_0332_ ;
 wire \u_ppwm/u_ex/_0333_ ;
 wire \u_ppwm/u_ex/_0334_ ;
 wire \u_ppwm/u_ex/_0335_ ;
 wire \u_ppwm/u_ex/_0336_ ;
 wire \u_ppwm/u_ex/_0337_ ;
 wire \u_ppwm/u_ex/_0338_ ;
 wire \u_ppwm/u_ex/_0339_ ;
 wire \u_ppwm/u_ex/_0340_ ;
 wire \u_ppwm/u_ex/_0341_ ;
 wire \u_ppwm/u_ex/_0342_ ;
 wire \u_ppwm/u_ex/_0343_ ;
 wire \u_ppwm/u_ex/_0344_ ;
 wire \u_ppwm/u_ex/_0345_ ;
 wire \u_ppwm/u_ex/_0346_ ;
 wire \u_ppwm/u_ex/_0347_ ;
 wire \u_ppwm/u_ex/_0348_ ;
 wire \u_ppwm/u_ex/_0349_ ;
 wire \u_ppwm/u_ex/_0350_ ;
 wire \u_ppwm/u_ex/_0351_ ;
 wire \u_ppwm/u_ex/_0352_ ;
 wire \u_ppwm/u_ex/_0353_ ;
 wire \u_ppwm/u_ex/_0354_ ;
 wire \u_ppwm/u_ex/_0355_ ;
 wire \u_ppwm/u_ex/_0356_ ;
 wire \u_ppwm/u_ex/_0357_ ;
 wire \u_ppwm/u_ex/_0358_ ;
 wire \u_ppwm/u_ex/_0359_ ;
 wire \u_ppwm/u_ex/_0360_ ;
 wire \u_ppwm/u_ex/_0361_ ;
 wire \u_ppwm/u_ex/_0362_ ;
 wire \u_ppwm/u_ex/_0363_ ;
 wire \u_ppwm/u_ex/_0364_ ;
 wire \u_ppwm/u_ex/_0365_ ;
 wire \u_ppwm/u_ex/_0366_ ;
 wire \u_ppwm/u_ex/_0367_ ;
 wire \u_ppwm/u_ex/_0368_ ;
 wire \u_ppwm/u_ex/_0369_ ;
 wire \u_ppwm/u_ex/_0370_ ;
 wire \u_ppwm/u_ex/_0371_ ;
 wire \u_ppwm/u_ex/_0372_ ;
 wire \u_ppwm/u_ex/_0373_ ;
 wire \u_ppwm/u_ex/_0374_ ;
 wire \u_ppwm/u_ex/_0375_ ;
 wire \u_ppwm/u_ex/_0376_ ;
 wire \u_ppwm/u_ex/_0377_ ;
 wire \u_ppwm/u_ex/_0378_ ;
 wire \u_ppwm/u_ex/_0379_ ;
 wire \u_ppwm/u_ex/_0380_ ;
 wire \u_ppwm/u_ex/_0381_ ;
 wire \u_ppwm/u_ex/_0382_ ;
 wire \u_ppwm/u_ex/_0383_ ;
 wire \u_ppwm/u_ex/_0384_ ;
 wire \u_ppwm/u_ex/_0385_ ;
 wire \u_ppwm/u_ex/_0386_ ;
 wire \u_ppwm/u_ex/_0387_ ;
 wire \u_ppwm/u_ex/_0388_ ;
 wire \u_ppwm/u_ex/_0389_ ;
 wire \u_ppwm/u_ex/_0390_ ;
 wire \u_ppwm/u_ex/_0391_ ;
 wire \u_ppwm/u_ex/_0392_ ;
 wire \u_ppwm/u_ex/_0393_ ;
 wire \u_ppwm/u_ex/_0394_ ;
 wire \u_ppwm/u_ex/_0395_ ;
 wire \u_ppwm/u_ex/_0396_ ;
 wire \u_ppwm/u_ex/_0397_ ;
 wire \u_ppwm/u_ex/_0398_ ;
 wire \u_ppwm/u_ex/_0399_ ;
 wire \u_ppwm/u_ex/_0400_ ;
 wire \u_ppwm/u_ex/_0401_ ;
 wire \u_ppwm/u_ex/_0402_ ;
 wire \u_ppwm/u_ex/_0403_ ;
 wire \u_ppwm/u_ex/_0404_ ;
 wire \u_ppwm/u_ex/_0405_ ;
 wire \u_ppwm/u_ex/_0406_ ;
 wire \u_ppwm/u_ex/_0407_ ;
 wire \u_ppwm/u_ex/_0408_ ;
 wire \u_ppwm/u_ex/_0409_ ;
 wire \u_ppwm/u_ex/_0410_ ;
 wire \u_ppwm/u_ex/_0411_ ;
 wire \u_ppwm/u_ex/_0412_ ;
 wire \u_ppwm/u_ex/_0413_ ;
 wire \u_ppwm/u_ex/_0414_ ;
 wire \u_ppwm/u_ex/_0415_ ;
 wire \u_ppwm/u_ex/_0416_ ;
 wire \u_ppwm/u_ex/_0417_ ;
 wire \u_ppwm/u_ex/_0418_ ;
 wire \u_ppwm/u_ex/_0419_ ;
 wire \u_ppwm/u_ex/_0420_ ;
 wire \u_ppwm/u_ex/_0421_ ;
 wire \u_ppwm/u_ex/_0422_ ;
 wire \u_ppwm/u_ex/_0423_ ;
 wire \u_ppwm/u_ex/_0424_ ;
 wire \u_ppwm/u_ex/_0425_ ;
 wire \u_ppwm/u_ex/_0426_ ;
 wire \u_ppwm/u_ex/_0427_ ;
 wire \u_ppwm/u_ex/_0428_ ;
 wire \u_ppwm/u_ex/_0429_ ;
 wire \u_ppwm/u_ex/_0430_ ;
 wire \u_ppwm/u_ex/_0431_ ;
 wire \u_ppwm/u_ex/_0432_ ;
 wire \u_ppwm/u_ex/_0433_ ;
 wire \u_ppwm/u_ex/_0434_ ;
 wire \u_ppwm/u_ex/_0435_ ;
 wire \u_ppwm/u_ex/_0436_ ;
 wire \u_ppwm/u_ex/_0437_ ;
 wire \u_ppwm/u_ex/_0438_ ;
 wire \u_ppwm/u_ex/_0439_ ;
 wire \u_ppwm/u_ex/_0440_ ;
 wire \u_ppwm/u_ex/_0441_ ;
 wire \u_ppwm/u_ex/_0442_ ;
 wire \u_ppwm/u_ex/_0443_ ;
 wire \u_ppwm/u_ex/_0444_ ;
 wire \u_ppwm/u_ex/_0445_ ;
 wire \u_ppwm/u_ex/_0446_ ;
 wire \u_ppwm/u_ex/_0447_ ;
 wire \u_ppwm/u_ex/_0448_ ;
 wire \u_ppwm/u_ex/_0449_ ;
 wire \u_ppwm/u_ex/_0450_ ;
 wire \u_ppwm/u_ex/_0451_ ;
 wire \u_ppwm/u_ex/_0452_ ;
 wire \u_ppwm/u_ex/_0453_ ;
 wire \u_ppwm/u_ex/_0454_ ;
 wire \u_ppwm/u_ex/_0455_ ;
 wire \u_ppwm/u_ex/_0456_ ;
 wire \u_ppwm/u_ex/_0457_ ;
 wire \u_ppwm/u_ex/_0458_ ;
 wire \u_ppwm/u_ex/_0459_ ;
 wire \u_ppwm/u_ex/_0460_ ;
 wire \u_ppwm/u_ex/_0461_ ;
 wire \u_ppwm/u_ex/_0462_ ;
 wire \u_ppwm/u_ex/_0463_ ;
 wire \u_ppwm/u_ex/_0464_ ;
 wire \u_ppwm/u_ex/_0465_ ;
 wire \u_ppwm/u_ex/_0466_ ;
 wire \u_ppwm/u_ex/_0467_ ;
 wire \u_ppwm/u_ex/_0468_ ;
 wire \u_ppwm/u_ex/_0469_ ;
 wire \u_ppwm/u_ex/_0470_ ;
 wire \u_ppwm/u_ex/_0471_ ;
 wire \u_ppwm/u_ex/_0472_ ;
 wire \u_ppwm/u_ex/_0473_ ;
 wire \u_ppwm/u_ex/_0474_ ;
 wire \u_ppwm/u_ex/_0475_ ;
 wire \u_ppwm/u_ex/_0476_ ;
 wire \u_ppwm/u_ex/_0477_ ;
 wire \u_ppwm/u_ex/_0478_ ;
 wire \u_ppwm/u_ex/_0479_ ;
 wire \u_ppwm/u_ex/_0480_ ;
 wire \u_ppwm/u_ex/_0481_ ;
 wire \u_ppwm/u_ex/_0482_ ;
 wire \u_ppwm/u_ex/_0483_ ;
 wire \u_ppwm/u_ex/_0484_ ;
 wire \u_ppwm/u_ex/_0485_ ;
 wire \u_ppwm/u_ex/_0486_ ;
 wire \u_ppwm/u_ex/_0487_ ;
 wire \u_ppwm/u_ex/_0488_ ;
 wire \u_ppwm/u_ex/_0489_ ;
 wire \u_ppwm/u_ex/_0490_ ;
 wire \u_ppwm/u_ex/_0491_ ;
 wire \u_ppwm/u_ex/_0492_ ;
 wire \u_ppwm/u_ex/_0493_ ;
 wire \u_ppwm/u_ex/_0494_ ;
 wire \u_ppwm/u_ex/_0495_ ;
 wire \u_ppwm/u_ex/_0496_ ;
 wire \u_ppwm/u_ex/_0497_ ;
 wire \u_ppwm/u_ex/_0498_ ;
 wire \u_ppwm/u_ex/_0499_ ;
 wire \u_ppwm/u_ex/_0500_ ;
 wire \u_ppwm/u_ex/_0501_ ;
 wire \u_ppwm/u_ex/_0502_ ;
 wire \u_ppwm/u_ex/_0503_ ;
 wire \u_ppwm/u_ex/_0504_ ;
 wire \u_ppwm/u_ex/_0505_ ;
 wire \u_ppwm/u_ex/_0506_ ;
 wire \u_ppwm/u_ex/_0507_ ;
 wire \u_ppwm/u_ex/_0508_ ;
 wire \u_ppwm/u_ex/_0509_ ;
 wire \u_ppwm/u_ex/_0510_ ;
 wire \u_ppwm/u_ex/_0511_ ;
 wire \u_ppwm/u_ex/_0512_ ;
 wire \u_ppwm/u_ex/_0513_ ;
 wire \u_ppwm/u_ex/_0514_ ;
 wire \u_ppwm/u_ex/_0515_ ;
 wire \u_ppwm/u_ex/_0516_ ;
 wire \u_ppwm/u_ex/_0517_ ;
 wire \u_ppwm/u_ex/_0518_ ;
 wire \u_ppwm/u_ex/_0519_ ;
 wire \u_ppwm/u_ex/_0520_ ;
 wire \u_ppwm/u_ex/_0521_ ;
 wire \u_ppwm/u_ex/_0522_ ;
 wire \u_ppwm/u_ex/_0523_ ;
 wire \u_ppwm/u_ex/_0524_ ;
 wire \u_ppwm/u_ex/_0525_ ;
 wire \u_ppwm/u_ex/_0526_ ;
 wire \u_ppwm/u_ex/_0527_ ;
 wire \u_ppwm/u_ex/_0528_ ;
 wire \u_ppwm/u_ex/_0529_ ;
 wire \u_ppwm/u_ex/_0530_ ;
 wire \u_ppwm/u_ex/_0531_ ;
 wire \u_ppwm/u_ex/_0532_ ;
 wire \u_ppwm/u_ex/_0533_ ;
 wire \u_ppwm/u_ex/_0534_ ;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire \u_ppwm/u_ex/cmp_flag_q ;
 wire \u_ppwm/u_ex/reg_value_q[0] ;
 wire \u_ppwm/u_ex/reg_value_q[1] ;
 wire \u_ppwm/u_ex/reg_value_q[2] ;
 wire \u_ppwm/u_ex/reg_value_q[3] ;
 wire \u_ppwm/u_ex/reg_value_q[4] ;
 wire \u_ppwm/u_ex/reg_value_q[5] ;
 wire \u_ppwm/u_ex/reg_value_q[6] ;
 wire \u_ppwm/u_ex/reg_value_q[7] ;
 wire \u_ppwm/u_ex/reg_value_q[8] ;
 wire \u_ppwm/u_ex/reg_value_q[9] ;
 wire \u_ppwm/u_ex/state_q[0] ;
 wire \u_ppwm/u_ex/state_q[1] ;
 wire \u_ppwm/u_ex/state_q[2] ;
 wire \u_ppwm/u_global_counter/_000_ ;
 wire \u_ppwm/u_global_counter/_001_ ;
 wire \u_ppwm/u_global_counter/_002_ ;
 wire \u_ppwm/u_global_counter/_003_ ;
 wire \u_ppwm/u_global_counter/_004_ ;
 wire \u_ppwm/u_global_counter/_005_ ;
 wire \u_ppwm/u_global_counter/_006_ ;
 wire \u_ppwm/u_global_counter/_007_ ;
 wire \u_ppwm/u_global_counter/_008_ ;
 wire \u_ppwm/u_global_counter/_009_ ;
 wire \u_ppwm/u_global_counter/_010_ ;
 wire \u_ppwm/u_global_counter/_011_ ;
 wire \u_ppwm/u_global_counter/_012_ ;
 wire \u_ppwm/u_global_counter/_013_ ;
 wire \u_ppwm/u_global_counter/_014_ ;
 wire \u_ppwm/u_global_counter/_015_ ;
 wire \u_ppwm/u_global_counter/_016_ ;
 wire \u_ppwm/u_global_counter/_017_ ;
 wire \u_ppwm/u_global_counter/_018_ ;
 wire \u_ppwm/u_global_counter/_019_ ;
 wire \u_ppwm/u_global_counter/_020_ ;
 wire \u_ppwm/u_global_counter/_021_ ;
 wire \u_ppwm/u_global_counter/_022_ ;
 wire \u_ppwm/u_global_counter/_023_ ;
 wire \u_ppwm/u_global_counter/_024_ ;
 wire \u_ppwm/u_global_counter/_025_ ;
 wire \u_ppwm/u_global_counter/_026_ ;
 wire \u_ppwm/u_global_counter/_027_ ;
 wire \u_ppwm/u_global_counter/_028_ ;
 wire \u_ppwm/u_global_counter/_029_ ;
 wire \u_ppwm/u_global_counter/_030_ ;
 wire \u_ppwm/u_global_counter/_031_ ;
 wire \u_ppwm/u_global_counter/_032_ ;
 wire \u_ppwm/u_global_counter/_033_ ;
 wire \u_ppwm/u_global_counter/_034_ ;
 wire \u_ppwm/u_global_counter/_035_ ;
 wire \u_ppwm/u_global_counter/_036_ ;
 wire \u_ppwm/u_global_counter/_037_ ;
 wire \u_ppwm/u_global_counter/_038_ ;
 wire \u_ppwm/u_global_counter/_039_ ;
 wire \u_ppwm/u_global_counter/_040_ ;
 wire \u_ppwm/u_global_counter/_041_ ;
 wire \u_ppwm/u_global_counter/_042_ ;
 wire \u_ppwm/u_global_counter/_043_ ;
 wire \u_ppwm/u_global_counter/_044_ ;
 wire \u_ppwm/u_global_counter/_045_ ;
 wire \u_ppwm/u_global_counter/_046_ ;
 wire \u_ppwm/u_global_counter/_047_ ;
 wire \u_ppwm/u_global_counter/_048_ ;
 wire \u_ppwm/u_global_counter/_049_ ;
 wire \u_ppwm/u_global_counter/_050_ ;
 wire \u_ppwm/u_global_counter/_051_ ;
 wire \u_ppwm/u_global_counter/_052_ ;
 wire \u_ppwm/u_mem/_0000_ ;
 wire \u_ppwm/u_mem/_0001_ ;
 wire \u_ppwm/u_mem/_0002_ ;
 wire \u_ppwm/u_mem/_0003_ ;
 wire \u_ppwm/u_mem/_0004_ ;
 wire \u_ppwm/u_mem/_0005_ ;
 wire \u_ppwm/u_mem/_0006_ ;
 wire \u_ppwm/u_mem/_0007_ ;
 wire \u_ppwm/u_mem/_0008_ ;
 wire \u_ppwm/u_mem/_0009_ ;
 wire \u_ppwm/u_mem/_0010_ ;
 wire \u_ppwm/u_mem/_0011_ ;
 wire \u_ppwm/u_mem/_0012_ ;
 wire \u_ppwm/u_mem/_0013_ ;
 wire \u_ppwm/u_mem/_0014_ ;
 wire \u_ppwm/u_mem/_0015_ ;
 wire \u_ppwm/u_mem/_0016_ ;
 wire \u_ppwm/u_mem/_0017_ ;
 wire \u_ppwm/u_mem/_0018_ ;
 wire \u_ppwm/u_mem/_0019_ ;
 wire \u_ppwm/u_mem/_0020_ ;
 wire \u_ppwm/u_mem/_0021_ ;
 wire \u_ppwm/u_mem/_0022_ ;
 wire \u_ppwm/u_mem/_0023_ ;
 wire \u_ppwm/u_mem/_0024_ ;
 wire \u_ppwm/u_mem/_0025_ ;
 wire \u_ppwm/u_mem/_0026_ ;
 wire \u_ppwm/u_mem/_0027_ ;
 wire \u_ppwm/u_mem/_0028_ ;
 wire \u_ppwm/u_mem/_0029_ ;
 wire \u_ppwm/u_mem/_0030_ ;
 wire \u_ppwm/u_mem/_0031_ ;
 wire \u_ppwm/u_mem/_0032_ ;
 wire \u_ppwm/u_mem/_0033_ ;
 wire \u_ppwm/u_mem/_0034_ ;
 wire \u_ppwm/u_mem/_0035_ ;
 wire \u_ppwm/u_mem/_0036_ ;
 wire \u_ppwm/u_mem/_0037_ ;
 wire \u_ppwm/u_mem/_0038_ ;
 wire \u_ppwm/u_mem/_0039_ ;
 wire \u_ppwm/u_mem/_0040_ ;
 wire \u_ppwm/u_mem/_0041_ ;
 wire \u_ppwm/u_mem/_0042_ ;
 wire \u_ppwm/u_mem/_0043_ ;
 wire \u_ppwm/u_mem/_0044_ ;
 wire \u_ppwm/u_mem/_0045_ ;
 wire \u_ppwm/u_mem/_0046_ ;
 wire \u_ppwm/u_mem/_0047_ ;
 wire \u_ppwm/u_mem/_0048_ ;
 wire \u_ppwm/u_mem/_0049_ ;
 wire \u_ppwm/u_mem/_0050_ ;
 wire \u_ppwm/u_mem/_0051_ ;
 wire \u_ppwm/u_mem/_0052_ ;
 wire \u_ppwm/u_mem/_0053_ ;
 wire \u_ppwm/u_mem/_0054_ ;
 wire \u_ppwm/u_mem/_0055_ ;
 wire \u_ppwm/u_mem/_0056_ ;
 wire \u_ppwm/u_mem/_0057_ ;
 wire \u_ppwm/u_mem/_0058_ ;
 wire \u_ppwm/u_mem/_0059_ ;
 wire \u_ppwm/u_mem/_0060_ ;
 wire \u_ppwm/u_mem/_0061_ ;
 wire \u_ppwm/u_mem/_0062_ ;
 wire \u_ppwm/u_mem/_0063_ ;
 wire \u_ppwm/u_mem/_0064_ ;
 wire \u_ppwm/u_mem/_0065_ ;
 wire \u_ppwm/u_mem/_0066_ ;
 wire \u_ppwm/u_mem/_0067_ ;
 wire \u_ppwm/u_mem/_0068_ ;
 wire \u_ppwm/u_mem/_0069_ ;
 wire \u_ppwm/u_mem/_0070_ ;
 wire \u_ppwm/u_mem/_0071_ ;
 wire \u_ppwm/u_mem/_0072_ ;
 wire \u_ppwm/u_mem/_0073_ ;
 wire \u_ppwm/u_mem/_0074_ ;
 wire \u_ppwm/u_mem/_0075_ ;
 wire \u_ppwm/u_mem/_0076_ ;
 wire \u_ppwm/u_mem/_0077_ ;
 wire \u_ppwm/u_mem/_0078_ ;
 wire \u_ppwm/u_mem/_0079_ ;
 wire \u_ppwm/u_mem/_0080_ ;
 wire \u_ppwm/u_mem/_0081_ ;
 wire \u_ppwm/u_mem/_0082_ ;
 wire \u_ppwm/u_mem/_0083_ ;
 wire \u_ppwm/u_mem/_0084_ ;
 wire \u_ppwm/u_mem/_0085_ ;
 wire \u_ppwm/u_mem/_0086_ ;
 wire \u_ppwm/u_mem/_0087_ ;
 wire \u_ppwm/u_mem/_0088_ ;
 wire \u_ppwm/u_mem/_0089_ ;
 wire \u_ppwm/u_mem/_0090_ ;
 wire \u_ppwm/u_mem/_0091_ ;
 wire \u_ppwm/u_mem/_0092_ ;
 wire \u_ppwm/u_mem/_0093_ ;
 wire \u_ppwm/u_mem/_0094_ ;
 wire \u_ppwm/u_mem/_0095_ ;
 wire \u_ppwm/u_mem/_0096_ ;
 wire \u_ppwm/u_mem/_0097_ ;
 wire \u_ppwm/u_mem/_0098_ ;
 wire \u_ppwm/u_mem/_0099_ ;
 wire \u_ppwm/u_mem/_0100_ ;
 wire \u_ppwm/u_mem/_0101_ ;
 wire \u_ppwm/u_mem/_0102_ ;
 wire \u_ppwm/u_mem/_0103_ ;
 wire \u_ppwm/u_mem/_0104_ ;
 wire \u_ppwm/u_mem/_0105_ ;
 wire \u_ppwm/u_mem/_0106_ ;
 wire \u_ppwm/u_mem/_0107_ ;
 wire \u_ppwm/u_mem/_0108_ ;
 wire \u_ppwm/u_mem/_0109_ ;
 wire \u_ppwm/u_mem/_0110_ ;
 wire \u_ppwm/u_mem/_0111_ ;
 wire \u_ppwm/u_mem/_0112_ ;
 wire \u_ppwm/u_mem/_0113_ ;
 wire \u_ppwm/u_mem/_0114_ ;
 wire \u_ppwm/u_mem/_0115_ ;
 wire \u_ppwm/u_mem/_0116_ ;
 wire \u_ppwm/u_mem/_0117_ ;
 wire \u_ppwm/u_mem/_0118_ ;
 wire \u_ppwm/u_mem/_0119_ ;
 wire \u_ppwm/u_mem/_0120_ ;
 wire \u_ppwm/u_mem/_0121_ ;
 wire \u_ppwm/u_mem/_0122_ ;
 wire \u_ppwm/u_mem/_0123_ ;
 wire \u_ppwm/u_mem/_0124_ ;
 wire \u_ppwm/u_mem/_0125_ ;
 wire \u_ppwm/u_mem/_0126_ ;
 wire \u_ppwm/u_mem/_0127_ ;
 wire \u_ppwm/u_mem/_0128_ ;
 wire \u_ppwm/u_mem/_0129_ ;
 wire \u_ppwm/u_mem/_0130_ ;
 wire \u_ppwm/u_mem/_0131_ ;
 wire \u_ppwm/u_mem/_0132_ ;
 wire \u_ppwm/u_mem/_0133_ ;
 wire \u_ppwm/u_mem/_0134_ ;
 wire \u_ppwm/u_mem/_0135_ ;
 wire \u_ppwm/u_mem/_0136_ ;
 wire \u_ppwm/u_mem/_0137_ ;
 wire \u_ppwm/u_mem/_0138_ ;
 wire \u_ppwm/u_mem/_0139_ ;
 wire \u_ppwm/u_mem/_0140_ ;
 wire \u_ppwm/u_mem/_0141_ ;
 wire \u_ppwm/u_mem/_0142_ ;
 wire \u_ppwm/u_mem/_0143_ ;
 wire \u_ppwm/u_mem/_0144_ ;
 wire \u_ppwm/u_mem/_0145_ ;
 wire \u_ppwm/u_mem/_0146_ ;
 wire \u_ppwm/u_mem/_0147_ ;
 wire \u_ppwm/u_mem/_0148_ ;
 wire \u_ppwm/u_mem/_0149_ ;
 wire \u_ppwm/u_mem/_0150_ ;
 wire \u_ppwm/u_mem/_0151_ ;
 wire \u_ppwm/u_mem/_0152_ ;
 wire \u_ppwm/u_mem/_0153_ ;
 wire \u_ppwm/u_mem/_0154_ ;
 wire \u_ppwm/u_mem/_0155_ ;
 wire \u_ppwm/u_mem/_0156_ ;
 wire \u_ppwm/u_mem/_0157_ ;
 wire \u_ppwm/u_mem/_0158_ ;
 wire \u_ppwm/u_mem/_0159_ ;
 wire \u_ppwm/u_mem/_0160_ ;
 wire \u_ppwm/u_mem/_0161_ ;
 wire \u_ppwm/u_mem/_0162_ ;
 wire \u_ppwm/u_mem/_0163_ ;
 wire \u_ppwm/u_mem/_0164_ ;
 wire \u_ppwm/u_mem/_0165_ ;
 wire \u_ppwm/u_mem/_0166_ ;
 wire \u_ppwm/u_mem/_0167_ ;
 wire \u_ppwm/u_mem/_0168_ ;
 wire \u_ppwm/u_mem/_0169_ ;
 wire \u_ppwm/u_mem/_0170_ ;
 wire \u_ppwm/u_mem/_0171_ ;
 wire \u_ppwm/u_mem/_0172_ ;
 wire \u_ppwm/u_mem/_0173_ ;
 wire \u_ppwm/u_mem/_0174_ ;
 wire \u_ppwm/u_mem/_0175_ ;
 wire \u_ppwm/u_mem/_0176_ ;
 wire \u_ppwm/u_mem/_0177_ ;
 wire \u_ppwm/u_mem/_0178_ ;
 wire \u_ppwm/u_mem/_0179_ ;
 wire \u_ppwm/u_mem/_0180_ ;
 wire \u_ppwm/u_mem/_0181_ ;
 wire \u_ppwm/u_mem/_0182_ ;
 wire \u_ppwm/u_mem/_0183_ ;
 wire \u_ppwm/u_mem/_0184_ ;
 wire \u_ppwm/u_mem/_0185_ ;
 wire \u_ppwm/u_mem/_0186_ ;
 wire \u_ppwm/u_mem/_0187_ ;
 wire \u_ppwm/u_mem/_0188_ ;
 wire \u_ppwm/u_mem/_0189_ ;
 wire \u_ppwm/u_mem/_0190_ ;
 wire \u_ppwm/u_mem/_0191_ ;
 wire \u_ppwm/u_mem/_0192_ ;
 wire \u_ppwm/u_mem/_0193_ ;
 wire \u_ppwm/u_mem/_0194_ ;
 wire \u_ppwm/u_mem/_0195_ ;
 wire \u_ppwm/u_mem/_0196_ ;
 wire \u_ppwm/u_mem/_0197_ ;
 wire \u_ppwm/u_mem/_0198_ ;
 wire \u_ppwm/u_mem/_0199_ ;
 wire \u_ppwm/u_mem/_0200_ ;
 wire \u_ppwm/u_mem/_0201_ ;
 wire \u_ppwm/u_mem/_0202_ ;
 wire \u_ppwm/u_mem/_0203_ ;
 wire \u_ppwm/u_mem/_0204_ ;
 wire \u_ppwm/u_mem/_0205_ ;
 wire \u_ppwm/u_mem/_0206_ ;
 wire \u_ppwm/u_mem/_0207_ ;
 wire \u_ppwm/u_mem/_0208_ ;
 wire \u_ppwm/u_mem/_0209_ ;
 wire \u_ppwm/u_mem/_0210_ ;
 wire \u_ppwm/u_mem/_0211_ ;
 wire \u_ppwm/u_mem/_0212_ ;
 wire \u_ppwm/u_mem/_0213_ ;
 wire \u_ppwm/u_mem/_0214_ ;
 wire \u_ppwm/u_mem/_0215_ ;
 wire \u_ppwm/u_mem/_0216_ ;
 wire \u_ppwm/u_mem/_0217_ ;
 wire \u_ppwm/u_mem/_0218_ ;
 wire \u_ppwm/u_mem/_0219_ ;
 wire \u_ppwm/u_mem/_0220_ ;
 wire \u_ppwm/u_mem/_0221_ ;
 wire \u_ppwm/u_mem/_0222_ ;
 wire \u_ppwm/u_mem/_0223_ ;
 wire \u_ppwm/u_mem/_0224_ ;
 wire \u_ppwm/u_mem/_0225_ ;
 wire \u_ppwm/u_mem/_0226_ ;
 wire \u_ppwm/u_mem/_0227_ ;
 wire \u_ppwm/u_mem/_0228_ ;
 wire \u_ppwm/u_mem/_0229_ ;
 wire \u_ppwm/u_mem/_0230_ ;
 wire \u_ppwm/u_mem/_0231_ ;
 wire \u_ppwm/u_mem/_0232_ ;
 wire \u_ppwm/u_mem/_0233_ ;
 wire \u_ppwm/u_mem/_0234_ ;
 wire \u_ppwm/u_mem/_0235_ ;
 wire \u_ppwm/u_mem/_0236_ ;
 wire \u_ppwm/u_mem/_0237_ ;
 wire \u_ppwm/u_mem/_0238_ ;
 wire \u_ppwm/u_mem/_0239_ ;
 wire \u_ppwm/u_mem/_0240_ ;
 wire \u_ppwm/u_mem/_0241_ ;
 wire \u_ppwm/u_mem/_0242_ ;
 wire \u_ppwm/u_mem/_0243_ ;
 wire \u_ppwm/u_mem/_0244_ ;
 wire \u_ppwm/u_mem/_0245_ ;
 wire \u_ppwm/u_mem/_0246_ ;
 wire \u_ppwm/u_mem/_0247_ ;
 wire \u_ppwm/u_mem/_0248_ ;
 wire \u_ppwm/u_mem/_0249_ ;
 wire \u_ppwm/u_mem/_0250_ ;
 wire \u_ppwm/u_mem/_0251_ ;
 wire \u_ppwm/u_mem/_0252_ ;
 wire \u_ppwm/u_mem/_0253_ ;
 wire \u_ppwm/u_mem/_0254_ ;
 wire \u_ppwm/u_mem/_0255_ ;
 wire \u_ppwm/u_mem/_0256_ ;
 wire \u_ppwm/u_mem/_0257_ ;
 wire \u_ppwm/u_mem/_0258_ ;
 wire \u_ppwm/u_mem/_0259_ ;
 wire \u_ppwm/u_mem/_0260_ ;
 wire \u_ppwm/u_mem/_0261_ ;
 wire \u_ppwm/u_mem/_0262_ ;
 wire \u_ppwm/u_mem/_0263_ ;
 wire \u_ppwm/u_mem/_0264_ ;
 wire \u_ppwm/u_mem/_0265_ ;
 wire \u_ppwm/u_mem/_0266_ ;
 wire \u_ppwm/u_mem/_0267_ ;
 wire \u_ppwm/u_mem/_0268_ ;
 wire \u_ppwm/u_mem/_0269_ ;
 wire \u_ppwm/u_mem/_0270_ ;
 wire \u_ppwm/u_mem/_0271_ ;
 wire \u_ppwm/u_mem/_0272_ ;
 wire \u_ppwm/u_mem/_0273_ ;
 wire \u_ppwm/u_mem/_0274_ ;
 wire \u_ppwm/u_mem/_0275_ ;
 wire \u_ppwm/u_mem/_0276_ ;
 wire \u_ppwm/u_mem/_0277_ ;
 wire \u_ppwm/u_mem/_0278_ ;
 wire \u_ppwm/u_mem/_0279_ ;
 wire \u_ppwm/u_mem/_0280_ ;
 wire \u_ppwm/u_mem/_0281_ ;
 wire \u_ppwm/u_mem/_0282_ ;
 wire \u_ppwm/u_mem/_0283_ ;
 wire \u_ppwm/u_mem/_0284_ ;
 wire \u_ppwm/u_mem/_0285_ ;
 wire \u_ppwm/u_mem/_0286_ ;
 wire \u_ppwm/u_mem/_0287_ ;
 wire \u_ppwm/u_mem/_0288_ ;
 wire \u_ppwm/u_mem/_0289_ ;
 wire \u_ppwm/u_mem/_0290_ ;
 wire \u_ppwm/u_mem/_0291_ ;
 wire \u_ppwm/u_mem/_0292_ ;
 wire \u_ppwm/u_mem/_0293_ ;
 wire \u_ppwm/u_mem/_0294_ ;
 wire \u_ppwm/u_mem/_0295_ ;
 wire \u_ppwm/u_mem/_0296_ ;
 wire \u_ppwm/u_mem/_0297_ ;
 wire \u_ppwm/u_mem/_0298_ ;
 wire \u_ppwm/u_mem/_0299_ ;
 wire \u_ppwm/u_mem/_0300_ ;
 wire \u_ppwm/u_mem/_0301_ ;
 wire \u_ppwm/u_mem/_0302_ ;
 wire \u_ppwm/u_mem/_0303_ ;
 wire \u_ppwm/u_mem/_0304_ ;
 wire \u_ppwm/u_mem/_0305_ ;
 wire \u_ppwm/u_mem/_0306_ ;
 wire \u_ppwm/u_mem/_0307_ ;
 wire \u_ppwm/u_mem/_0308_ ;
 wire \u_ppwm/u_mem/_0309_ ;
 wire \u_ppwm/u_mem/_0310_ ;
 wire \u_ppwm/u_mem/_0311_ ;
 wire \u_ppwm/u_mem/_0312_ ;
 wire \u_ppwm/u_mem/_0313_ ;
 wire \u_ppwm/u_mem/_0314_ ;
 wire \u_ppwm/u_mem/_0315_ ;
 wire \u_ppwm/u_mem/_0316_ ;
 wire \u_ppwm/u_mem/_0317_ ;
 wire \u_ppwm/u_mem/_0318_ ;
 wire \u_ppwm/u_mem/_0319_ ;
 wire \u_ppwm/u_mem/_0320_ ;
 wire \u_ppwm/u_mem/_0321_ ;
 wire \u_ppwm/u_mem/_0322_ ;
 wire \u_ppwm/u_mem/_0323_ ;
 wire \u_ppwm/u_mem/_0324_ ;
 wire \u_ppwm/u_mem/_0325_ ;
 wire \u_ppwm/u_mem/_0326_ ;
 wire \u_ppwm/u_mem/_0327_ ;
 wire \u_ppwm/u_mem/_0328_ ;
 wire \u_ppwm/u_mem/_0329_ ;
 wire \u_ppwm/u_mem/_0330_ ;
 wire \u_ppwm/u_mem/_0331_ ;
 wire \u_ppwm/u_mem/_0332_ ;
 wire \u_ppwm/u_mem/_0333_ ;
 wire \u_ppwm/u_mem/_0334_ ;
 wire \u_ppwm/u_mem/_0335_ ;
 wire \u_ppwm/u_mem/_0336_ ;
 wire \u_ppwm/u_mem/_0337_ ;
 wire \u_ppwm/u_mem/_0338_ ;
 wire \u_ppwm/u_mem/_0339_ ;
 wire \u_ppwm/u_mem/_0340_ ;
 wire \u_ppwm/u_mem/_0341_ ;
 wire \u_ppwm/u_mem/_0342_ ;
 wire \u_ppwm/u_mem/_0343_ ;
 wire \u_ppwm/u_mem/_0344_ ;
 wire \u_ppwm/u_mem/_0345_ ;
 wire \u_ppwm/u_mem/_0346_ ;
 wire \u_ppwm/u_mem/_0347_ ;
 wire \u_ppwm/u_mem/_0348_ ;
 wire \u_ppwm/u_mem/_0349_ ;
 wire \u_ppwm/u_mem/_0350_ ;
 wire \u_ppwm/u_mem/_0351_ ;
 wire \u_ppwm/u_mem/_0352_ ;
 wire \u_ppwm/u_mem/_0353_ ;
 wire \u_ppwm/u_mem/_0354_ ;
 wire \u_ppwm/u_mem/_0355_ ;
 wire \u_ppwm/u_mem/_0356_ ;
 wire \u_ppwm/u_mem/_0357_ ;
 wire \u_ppwm/u_mem/_0358_ ;
 wire \u_ppwm/u_mem/_0359_ ;
 wire \u_ppwm/u_mem/_0360_ ;
 wire \u_ppwm/u_mem/_0361_ ;
 wire \u_ppwm/u_mem/_0362_ ;
 wire \u_ppwm/u_mem/_0363_ ;
 wire \u_ppwm/u_mem/_0364_ ;
 wire \u_ppwm/u_mem/_0365_ ;
 wire \u_ppwm/u_mem/_0366_ ;
 wire \u_ppwm/u_mem/_0367_ ;
 wire \u_ppwm/u_mem/_0368_ ;
 wire \u_ppwm/u_mem/_0369_ ;
 wire \u_ppwm/u_mem/_0370_ ;
 wire \u_ppwm/u_mem/_0371_ ;
 wire \u_ppwm/u_mem/_0372_ ;
 wire \u_ppwm/u_mem/_0373_ ;
 wire \u_ppwm/u_mem/_0374_ ;
 wire \u_ppwm/u_mem/_0375_ ;
 wire \u_ppwm/u_mem/_0376_ ;
 wire \u_ppwm/u_mem/_0377_ ;
 wire \u_ppwm/u_mem/_0378_ ;
 wire \u_ppwm/u_mem/_0379_ ;
 wire \u_ppwm/u_mem/_0380_ ;
 wire \u_ppwm/u_mem/_0381_ ;
 wire \u_ppwm/u_mem/_0382_ ;
 wire \u_ppwm/u_mem/_0383_ ;
 wire \u_ppwm/u_mem/_0384_ ;
 wire \u_ppwm/u_mem/_0385_ ;
 wire \u_ppwm/u_mem/_0386_ ;
 wire \u_ppwm/u_mem/_0387_ ;
 wire \u_ppwm/u_mem/_0388_ ;
 wire \u_ppwm/u_mem/_0389_ ;
 wire \u_ppwm/u_mem/_0390_ ;
 wire \u_ppwm/u_mem/_0391_ ;
 wire \u_ppwm/u_mem/_0392_ ;
 wire \u_ppwm/u_mem/_0393_ ;
 wire \u_ppwm/u_mem/_0394_ ;
 wire \u_ppwm/u_mem/_0395_ ;
 wire \u_ppwm/u_mem/_0396_ ;
 wire \u_ppwm/u_mem/_0397_ ;
 wire \u_ppwm/u_mem/_0398_ ;
 wire \u_ppwm/u_mem/_0399_ ;
 wire \u_ppwm/u_mem/_0400_ ;
 wire \u_ppwm/u_mem/_0401_ ;
 wire \u_ppwm/u_mem/_0402_ ;
 wire \u_ppwm/u_mem/_0403_ ;
 wire \u_ppwm/u_mem/_0404_ ;
 wire \u_ppwm/u_mem/_0405_ ;
 wire \u_ppwm/u_mem/_0406_ ;
 wire \u_ppwm/u_mem/_0407_ ;
 wire \u_ppwm/u_mem/_0408_ ;
 wire \u_ppwm/u_mem/_0409_ ;
 wire \u_ppwm/u_mem/_0410_ ;
 wire \u_ppwm/u_mem/_0411_ ;
 wire \u_ppwm/u_mem/_0412_ ;
 wire \u_ppwm/u_mem/_0413_ ;
 wire \u_ppwm/u_mem/_0414_ ;
 wire \u_ppwm/u_mem/_0415_ ;
 wire \u_ppwm/u_mem/_0416_ ;
 wire \u_ppwm/u_mem/_0417_ ;
 wire \u_ppwm/u_mem/_0418_ ;
 wire \u_ppwm/u_mem/_0419_ ;
 wire \u_ppwm/u_mem/_0420_ ;
 wire \u_ppwm/u_mem/_0421_ ;
 wire \u_ppwm/u_mem/_0422_ ;
 wire \u_ppwm/u_mem/_0423_ ;
 wire \u_ppwm/u_mem/_0424_ ;
 wire \u_ppwm/u_mem/_0425_ ;
 wire \u_ppwm/u_mem/_0426_ ;
 wire \u_ppwm/u_mem/_0427_ ;
 wire \u_ppwm/u_mem/_0428_ ;
 wire \u_ppwm/u_mem/_0429_ ;
 wire \u_ppwm/u_mem/_0430_ ;
 wire \u_ppwm/u_mem/_0431_ ;
 wire \u_ppwm/u_mem/_0432_ ;
 wire \u_ppwm/u_mem/_0433_ ;
 wire \u_ppwm/u_mem/_0434_ ;
 wire \u_ppwm/u_mem/_0435_ ;
 wire \u_ppwm/u_mem/_0436_ ;
 wire \u_ppwm/u_mem/_0437_ ;
 wire \u_ppwm/u_mem/_0438_ ;
 wire \u_ppwm/u_mem/_0439_ ;
 wire \u_ppwm/u_mem/_0440_ ;
 wire \u_ppwm/u_mem/_0441_ ;
 wire \u_ppwm/u_mem/_0442_ ;
 wire \u_ppwm/u_mem/_0443_ ;
 wire \u_ppwm/u_mem/_0444_ ;
 wire \u_ppwm/u_mem/_0445_ ;
 wire \u_ppwm/u_mem/_0446_ ;
 wire \u_ppwm/u_mem/_0447_ ;
 wire \u_ppwm/u_mem/_0448_ ;
 wire \u_ppwm/u_mem/_0449_ ;
 wire \u_ppwm/u_mem/_0450_ ;
 wire \u_ppwm/u_mem/_0451_ ;
 wire \u_ppwm/u_mem/_0452_ ;
 wire \u_ppwm/u_mem/_0453_ ;
 wire \u_ppwm/u_mem/_0454_ ;
 wire \u_ppwm/u_mem/_0455_ ;
 wire \u_ppwm/u_mem/_0456_ ;
 wire \u_ppwm/u_mem/_0457_ ;
 wire \u_ppwm/u_mem/_0458_ ;
 wire \u_ppwm/u_mem/_0459_ ;
 wire \u_ppwm/u_mem/_0460_ ;
 wire \u_ppwm/u_mem/_0461_ ;
 wire \u_ppwm/u_mem/_0462_ ;
 wire \u_ppwm/u_mem/_0463_ ;
 wire \u_ppwm/u_mem/_0464_ ;
 wire \u_ppwm/u_mem/_0465_ ;
 wire \u_ppwm/u_mem/_0466_ ;
 wire \u_ppwm/u_mem/_0467_ ;
 wire \u_ppwm/u_mem/_0468_ ;
 wire \u_ppwm/u_mem/_0469_ ;
 wire \u_ppwm/u_mem/_0470_ ;
 wire \u_ppwm/u_mem/_0471_ ;
 wire \u_ppwm/u_mem/_0472_ ;
 wire \u_ppwm/u_mem/_0473_ ;
 wire \u_ppwm/u_mem/_0474_ ;
 wire \u_ppwm/u_mem/_0475_ ;
 wire \u_ppwm/u_mem/_0476_ ;
 wire \u_ppwm/u_mem/_0477_ ;
 wire \u_ppwm/u_mem/_0478_ ;
 wire \u_ppwm/u_mem/_0479_ ;
 wire \u_ppwm/u_mem/_0480_ ;
 wire \u_ppwm/u_mem/_0481_ ;
 wire \u_ppwm/u_mem/_0482_ ;
 wire \u_ppwm/u_mem/_0483_ ;
 wire \u_ppwm/u_mem/_0484_ ;
 wire \u_ppwm/u_mem/_0485_ ;
 wire \u_ppwm/u_mem/_0486_ ;
 wire \u_ppwm/u_mem/_0487_ ;
 wire \u_ppwm/u_mem/_0488_ ;
 wire \u_ppwm/u_mem/_0489_ ;
 wire \u_ppwm/u_mem/_0490_ ;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire \u_ppwm/u_mem/bit_count[0] ;
 wire \u_ppwm/u_mem/bit_count[1] ;
 wire \u_ppwm/u_mem/bit_count[2] ;
 wire \u_ppwm/u_mem/bit_count[3] ;
 wire \u_ppwm/u_mem/bit_count[4] ;
 wire \u_ppwm/u_mem/bit_count[5] ;
 wire \u_ppwm/u_mem/bit_count[6] ;
 wire \u_ppwm/u_mem/memory[0] ;
 wire \u_ppwm/u_mem/memory[100] ;
 wire \u_ppwm/u_mem/memory[101] ;
 wire \u_ppwm/u_mem/memory[102] ;
 wire \u_ppwm/u_mem/memory[103] ;
 wire \u_ppwm/u_mem/memory[104] ;
 wire \u_ppwm/u_mem/memory[105] ;
 wire \u_ppwm/u_mem/memory[106] ;
 wire \u_ppwm/u_mem/memory[107] ;
 wire \u_ppwm/u_mem/memory[10] ;
 wire \u_ppwm/u_mem/memory[11] ;
 wire \u_ppwm/u_mem/memory[12] ;
 wire \u_ppwm/u_mem/memory[13] ;
 wire \u_ppwm/u_mem/memory[14] ;
 wire \u_ppwm/u_mem/memory[15] ;
 wire \u_ppwm/u_mem/memory[16] ;
 wire \u_ppwm/u_mem/memory[17] ;
 wire \u_ppwm/u_mem/memory[18] ;
 wire \u_ppwm/u_mem/memory[19] ;
 wire \u_ppwm/u_mem/memory[1] ;
 wire \u_ppwm/u_mem/memory[20] ;
 wire \u_ppwm/u_mem/memory[21] ;
 wire \u_ppwm/u_mem/memory[22] ;
 wire \u_ppwm/u_mem/memory[23] ;
 wire \u_ppwm/u_mem/memory[24] ;
 wire \u_ppwm/u_mem/memory[25] ;
 wire \u_ppwm/u_mem/memory[26] ;
 wire \u_ppwm/u_mem/memory[27] ;
 wire \u_ppwm/u_mem/memory[28] ;
 wire \u_ppwm/u_mem/memory[29] ;
 wire \u_ppwm/u_mem/memory[2] ;
 wire \u_ppwm/u_mem/memory[30] ;
 wire \u_ppwm/u_mem/memory[31] ;
 wire \u_ppwm/u_mem/memory[32] ;
 wire \u_ppwm/u_mem/memory[33] ;
 wire \u_ppwm/u_mem/memory[34] ;
 wire \u_ppwm/u_mem/memory[35] ;
 wire \u_ppwm/u_mem/memory[36] ;
 wire \u_ppwm/u_mem/memory[37] ;
 wire \u_ppwm/u_mem/memory[38] ;
 wire \u_ppwm/u_mem/memory[39] ;
 wire \u_ppwm/u_mem/memory[3] ;
 wire \u_ppwm/u_mem/memory[40] ;
 wire \u_ppwm/u_mem/memory[41] ;
 wire \u_ppwm/u_mem/memory[42] ;
 wire \u_ppwm/u_mem/memory[43] ;
 wire \u_ppwm/u_mem/memory[44] ;
 wire \u_ppwm/u_mem/memory[45] ;
 wire \u_ppwm/u_mem/memory[46] ;
 wire \u_ppwm/u_mem/memory[47] ;
 wire \u_ppwm/u_mem/memory[48] ;
 wire \u_ppwm/u_mem/memory[49] ;
 wire \u_ppwm/u_mem/memory[4] ;
 wire \u_ppwm/u_mem/memory[50] ;
 wire \u_ppwm/u_mem/memory[51] ;
 wire \u_ppwm/u_mem/memory[52] ;
 wire \u_ppwm/u_mem/memory[53] ;
 wire \u_ppwm/u_mem/memory[54] ;
 wire \u_ppwm/u_mem/memory[55] ;
 wire \u_ppwm/u_mem/memory[56] ;
 wire \u_ppwm/u_mem/memory[57] ;
 wire \u_ppwm/u_mem/memory[58] ;
 wire \u_ppwm/u_mem/memory[59] ;
 wire \u_ppwm/u_mem/memory[5] ;
 wire \u_ppwm/u_mem/memory[60] ;
 wire \u_ppwm/u_mem/memory[61] ;
 wire \u_ppwm/u_mem/memory[62] ;
 wire \u_ppwm/u_mem/memory[63] ;
 wire \u_ppwm/u_mem/memory[64] ;
 wire \u_ppwm/u_mem/memory[65] ;
 wire \u_ppwm/u_mem/memory[66] ;
 wire \u_ppwm/u_mem/memory[67] ;
 wire \u_ppwm/u_mem/memory[68] ;
 wire \u_ppwm/u_mem/memory[69] ;
 wire \u_ppwm/u_mem/memory[6] ;
 wire \u_ppwm/u_mem/memory[70] ;
 wire \u_ppwm/u_mem/memory[71] ;
 wire \u_ppwm/u_mem/memory[72] ;
 wire \u_ppwm/u_mem/memory[73] ;
 wire \u_ppwm/u_mem/memory[74] ;
 wire \u_ppwm/u_mem/memory[75] ;
 wire \u_ppwm/u_mem/memory[76] ;
 wire \u_ppwm/u_mem/memory[77] ;
 wire \u_ppwm/u_mem/memory[78] ;
 wire \u_ppwm/u_mem/memory[79] ;
 wire \u_ppwm/u_mem/memory[7] ;
 wire \u_ppwm/u_mem/memory[80] ;
 wire \u_ppwm/u_mem/memory[81] ;
 wire \u_ppwm/u_mem/memory[82] ;
 wire \u_ppwm/u_mem/memory[83] ;
 wire \u_ppwm/u_mem/memory[84] ;
 wire \u_ppwm/u_mem/memory[85] ;
 wire \u_ppwm/u_mem/memory[86] ;
 wire \u_ppwm/u_mem/memory[87] ;
 wire \u_ppwm/u_mem/memory[88] ;
 wire \u_ppwm/u_mem/memory[89] ;
 wire \u_ppwm/u_mem/memory[8] ;
 wire \u_ppwm/u_mem/memory[90] ;
 wire \u_ppwm/u_mem/memory[91] ;
 wire \u_ppwm/u_mem/memory[92] ;
 wire \u_ppwm/u_mem/memory[93] ;
 wire \u_ppwm/u_mem/memory[94] ;
 wire \u_ppwm/u_mem/memory[95] ;
 wire \u_ppwm/u_mem/memory[96] ;
 wire \u_ppwm/u_mem/memory[97] ;
 wire \u_ppwm/u_mem/memory[98] ;
 wire \u_ppwm/u_mem/memory[99] ;
 wire \u_ppwm/u_mem/memory[9] ;
 wire \u_ppwm/u_mem/state_q[0] ;
 wire \u_ppwm/u_mem/state_q[2] ;
 wire \u_ppwm/u_pwm/_000_ ;
 wire \u_ppwm/u_pwm/_001_ ;
 wire \u_ppwm/u_pwm/_002_ ;
 wire \u_ppwm/u_pwm/_003_ ;
 wire \u_ppwm/u_pwm/_004_ ;
 wire \u_ppwm/u_pwm/_005_ ;
 wire \u_ppwm/u_pwm/_006_ ;
 wire \u_ppwm/u_pwm/_007_ ;
 wire \u_ppwm/u_pwm/_008_ ;
 wire \u_ppwm/u_pwm/_009_ ;
 wire \u_ppwm/u_pwm/_010_ ;
 wire \u_ppwm/u_pwm/_011_ ;
 wire \u_ppwm/u_pwm/_012_ ;
 wire \u_ppwm/u_pwm/_013_ ;
 wire \u_ppwm/u_pwm/_014_ ;
 wire \u_ppwm/u_pwm/_015_ ;
 wire \u_ppwm/u_pwm/_016_ ;
 wire \u_ppwm/u_pwm/_017_ ;
 wire \u_ppwm/u_pwm/_018_ ;
 wire \u_ppwm/u_pwm/_019_ ;
 wire \u_ppwm/u_pwm/_020_ ;
 wire \u_ppwm/u_pwm/_021_ ;
 wire \u_ppwm/u_pwm/_022_ ;
 wire \u_ppwm/u_pwm/_023_ ;
 wire \u_ppwm/u_pwm/_024_ ;
 wire \u_ppwm/u_pwm/_025_ ;
 wire \u_ppwm/u_pwm/_026_ ;
 wire \u_ppwm/u_pwm/_027_ ;
 wire \u_ppwm/u_pwm/_028_ ;
 wire \u_ppwm/u_pwm/_029_ ;
 wire \u_ppwm/u_pwm/_030_ ;
 wire \u_ppwm/u_pwm/_031_ ;
 wire \u_ppwm/u_pwm/_032_ ;
 wire \u_ppwm/u_pwm/_033_ ;
 wire \u_ppwm/u_pwm/_034_ ;
 wire \u_ppwm/u_pwm/_035_ ;
 wire \u_ppwm/u_pwm/_036_ ;
 wire \u_ppwm/u_pwm/_037_ ;
 wire \u_ppwm/u_pwm/_038_ ;
 wire \u_ppwm/u_pwm/_039_ ;
 wire \u_ppwm/u_pwm/_040_ ;
 wire \u_ppwm/u_pwm/_041_ ;
 wire \u_ppwm/u_pwm/_042_ ;
 wire \u_ppwm/u_pwm/_043_ ;
 wire \u_ppwm/u_pwm/_044_ ;
 wire \u_ppwm/u_pwm/_045_ ;
 wire \u_ppwm/u_pwm/_046_ ;
 wire \u_ppwm/u_pwm/_047_ ;
 wire \u_ppwm/u_pwm/_048_ ;
 wire \u_ppwm/u_pwm/_049_ ;
 wire \u_ppwm/u_pwm/_050_ ;
 wire \u_ppwm/u_pwm/_051_ ;
 wire \u_ppwm/u_pwm/_052_ ;
 wire \u_ppwm/u_pwm/_053_ ;
 wire \u_ppwm/u_pwm/_054_ ;
 wire \u_ppwm/u_pwm/_055_ ;
 wire \u_ppwm/u_pwm/_056_ ;
 wire \u_ppwm/u_pwm/_057_ ;
 wire \u_ppwm/u_pwm/_058_ ;
 wire \u_ppwm/u_pwm/_059_ ;
 wire \u_ppwm/u_pwm/_060_ ;
 wire \u_ppwm/u_pwm/_061_ ;
 wire \u_ppwm/u_pwm/_062_ ;
 wire \u_ppwm/u_pwm/_063_ ;
 wire \u_ppwm/u_pwm/_064_ ;
 wire \u_ppwm/u_pwm/_065_ ;
 wire \u_ppwm/u_pwm/_066_ ;
 wire \u_ppwm/u_pwm/_067_ ;
 wire \u_ppwm/u_pwm/_068_ ;
 wire \u_ppwm/u_pwm/_069_ ;
 wire \u_ppwm/u_pwm/_070_ ;
 wire \u_ppwm/u_pwm/_071_ ;
 wire \u_ppwm/u_pwm/_072_ ;
 wire \u_ppwm/u_pwm/_073_ ;
 wire \u_ppwm/u_pwm/_074_ ;
 wire \u_ppwm/u_pwm/_075_ ;
 wire \u_ppwm/u_pwm/_076_ ;
 wire \u_ppwm/u_pwm/_077_ ;
 wire \u_ppwm/u_pwm/_078_ ;
 wire \u_ppwm/u_pwm/_079_ ;
 wire \u_ppwm/u_pwm/_080_ ;
 wire \u_ppwm/u_pwm/_081_ ;
 wire \u_ppwm/u_pwm/_082_ ;
 wire \u_ppwm/u_pwm/_083_ ;
 wire \u_ppwm/u_pwm/_084_ ;
 wire \u_ppwm/u_pwm/_085_ ;
 wire \u_ppwm/u_pwm/_086_ ;
 wire \u_ppwm/u_pwm/_087_ ;
 wire \u_ppwm/u_pwm/_088_ ;
 wire \u_ppwm/u_pwm/_089_ ;
 wire \u_ppwm/u_pwm/_090_ ;
 wire \u_ppwm/u_pwm/_091_ ;
 wire \u_ppwm/u_pwm/_092_ ;
 wire \u_ppwm/u_pwm/_093_ ;
 wire \u_ppwm/u_pwm/_094_ ;
 wire \u_ppwm/u_pwm/_095_ ;
 wire \u_ppwm/u_pwm/_096_ ;
 wire \u_ppwm/u_pwm/_097_ ;
 wire \u_ppwm/u_pwm/_098_ ;
 wire \u_ppwm/u_pwm/_099_ ;
 wire \u_ppwm/u_pwm/_100_ ;
 wire \u_ppwm/u_pwm/_101_ ;
 wire \u_ppwm/u_pwm/_102_ ;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire clknet_0_clk;
 wire \u_ppwm/u_pwm/cmp_value[0] ;
 wire \u_ppwm/u_pwm/cmp_value[1] ;
 wire \u_ppwm/u_pwm/cmp_value[2] ;
 wire \u_ppwm/u_pwm/cmp_value[3] ;
 wire \u_ppwm/u_pwm/cmp_value[4] ;
 wire \u_ppwm/u_pwm/cmp_value[5] ;
 wire \u_ppwm/u_pwm/cmp_value[6] ;
 wire \u_ppwm/u_pwm/cmp_value[7] ;
 wire \u_ppwm/u_pwm/cmp_value[8] ;
 wire \u_ppwm/u_pwm/cmp_value[9] ;
 wire \u_ppwm/u_pwm/counter[0] ;
 wire \u_ppwm/u_pwm/counter[1] ;
 wire \u_ppwm/u_pwm/counter[2] ;
 wire \u_ppwm/u_pwm/counter[3] ;
 wire \u_ppwm/u_pwm/counter[4] ;
 wire \u_ppwm/u_pwm/counter[5] ;
 wire \u_ppwm/u_pwm/counter[6] ;
 wire \u_ppwm/u_pwm/counter[7] ;
 wire \u_ppwm/u_pwm/counter[8] ;
 wire \u_ppwm/u_pwm/counter[9] ;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net1;
 wire net3;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;

 sg13g2_tielo heichips25_ppwm_4 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net4));
 sg13g2_tielo heichips25_ppwm_5 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net5));
 sg13g2_tielo heichips25_ppwm_6 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net6));
 sg13g2_tielo heichips25_ppwm_7 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net7));
 sg13g2_tielo heichips25_ppwm_8 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net8));
 sg13g2_tielo heichips25_ppwm_9 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net9));
 sg13g2_tielo heichips25_ppwm_10 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net10));
 sg13g2_tielo heichips25_ppwm_11 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net11));
 sg13g2_tielo heichips25_ppwm_12 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net12));
 sg13g2_tielo heichips25_ppwm_13 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net13));
 sg13g2_tielo heichips25_ppwm_14 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net14));
 sg13g2_tielo heichips25_ppwm_15 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net15));
 sg13g2_tielo heichips25_ppwm_16 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net16));
 sg13g2_tielo heichips25_ppwm_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net17));
 sg13g2_tielo heichips25_ppwm_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net18));
 sg13g2_tielo heichips25_ppwm_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net19));
 sg13g2_tielo heichips25_ppwm_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net20));
 sg13g2_tielo heichips25_ppwm_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net21));
 sg13g2_tielo heichips25_ppwm_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net22));
 sg13g2_tielo heichips25_ppwm_23 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net23));
 sg13g2_tielo heichips25_ppwm_24 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net24));
 sg13g2_tielo heichips25_ppwm_25 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net25));
 sg13g2_tiehi \u_ppwm/u_ex/_1119__26  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net26));
 sg13g2_inv_2 \u_ppwm/u_ex/_0564_  (.Y(\u_ppwm/u_ex/_0523_ ),
    .A(\u_ppwm/u_ex/reg_value_q[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_ex/_0565_  (.Y(\u_ppwm/u_ex/_0524_ ),
    .A(\u_ppwm/u_ex/reg_value_q[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 \u_ppwm/u_ex/_0566_  (.A(\u_ppwm/u_ex/reg_value_q[7] ),
    .Y(\u_ppwm/u_ex/_0525_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_ex/_0567_  (.Y(\u_ppwm/u_ex/_0526_ ),
    .A(net448),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 \u_ppwm/u_ex/_0568_  (.A(\u_ppwm/u_ex/reg_value_q[5] ),
    .Y(\u_ppwm/u_ex/_0527_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_ex/_0569_  (.Y(\u_ppwm/u_ex/_0528_ ),
    .A(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0570_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0529_ ),
    .A(net451),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0571_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0530_ ),
    .A(net454),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_ex/_0572_  (.Y(\u_ppwm/u_ex/_0531_ ),
    .A(net455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_ex/_0573_  (.Y(\u_ppwm/u_ex/_0532_ ),
    .A(\u_ppwm/pwm_value[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0574_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0533_ ),
    .A(net458),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0575_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0534_ ),
    .A(net460),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0576_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0029_ ),
    .A(net462),
    .VSS(VGND));
 sg13g2_inv_4 \u_ppwm/u_ex/_0577_  (.A(net463),
    .Y(\u_ppwm/u_ex/_0030_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0578_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0031_ ),
    .A(net247),
    .VSS(VGND));
 sg13g2_inv_4 \u_ppwm/u_ex/_0579_  (.A(net506),
    .Y(\u_ppwm/u_ex/_0032_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0580_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0033_ ),
    .A(\u_ppwm/instr[0] ),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_ex/_0581_  (.Y(\u_ppwm/u_ex/_0034_ ),
    .A(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 \u_ppwm/u_ex/_0582_  (.A(net373),
    .Y(\u_ppwm/u_ex/_0035_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0583_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0036_ ),
    .A(net377),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0584_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0037_ ),
    .A(net399),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0585_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0038_ ),
    .A(\u_ppwm/global_counter[18] ),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0586_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0039_ ),
    .A(\u_ppwm/global_counter[14] ),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0587_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0040_ ),
    .A(net440),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0588_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0041_ ),
    .A(\u_ppwm/global_counter[6] ),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0589_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0042_ ),
    .A(\u_ppwm/global_counter[4] ),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0590_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0043_ ),
    .A(\u_ppwm/global_counter[3] ),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0591_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0044_ ),
    .A(net443),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0592_  (.B1(net399),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0045_ ),
    .VSS(VGND),
    .A1(net217),
    .A2(net614));
 sg13g2_and2_1 \u_ppwm/u_ex/_0593_  (.A(net473),
    .B(net480),
    .X(\u_ppwm/u_ex/_0046_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_ex/_0594_  (.B(net469),
    .C(\u_ppwm/u_ex/_0046_ ),
    .A(net468),
    .Y(\u_ppwm/u_ex/_0047_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 \u_ppwm/u_ex/_0595_  (.A(\u_ppwm/instr[0] ),
    .B(\u_ppwm/instr[1] ),
    .Y(\u_ppwm/u_ex/_0048_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0596_  (.A(net388),
    .B(\u_ppwm/instr[0] ),
    .C(\u_ppwm/instr[1] ),
    .Y(\u_ppwm/u_ex/_0049_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 \u_ppwm/u_ex/_0597_  (.A(net381),
    .B_N(net384),
    .Y(\u_ppwm/u_ex/_0050_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0598_  (.A(net375),
    .B(net378),
    .Y(\u_ppwm/u_ex/_0051_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_ex/_0599_  (.B(\u_ppwm/u_ex/_0050_ ),
    .C(net369),
    .A(\u_ppwm/u_ex/_0049_ ),
    .Y(\u_ppwm/u_ex/_0052_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0600_  (.Y(\u_ppwm/u_ex/_0053_ ),
    .A(net446),
    .B(\u_ppwm/u_ex/_0052_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_ex/_0601_  (.B(\u_ppwm/u_ex/_0047_ ),
    .C(\u_ppwm/u_ex/_0052_ ),
    .A(net446),
    .Y(\u_ppwm/u_ex/_0054_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0602_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0045_ ),
    .A2(\u_ppwm/u_ex/_0054_ ),
    .Y(\u_ppwm/u_ex/_0002_ ),
    .B1(\u_ppwm/u_ex/_0032_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0603_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0037_ ),
    .A2(net614),
    .Y(\u_ppwm/u_ex/_0055_ ),
    .B1(\u_ppwm/u_ex/_0032_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0604_  (.B1(net615),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0000_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0047_ ),
    .A2(\u_ppwm/u_ex/_0053_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0605_  (.Y(\u_ppwm/u_ex/_0056_ ),
    .A(\u_ppwm/u_ex/_0037_ ),
    .B(net217),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_ex/_0606_  (.B(\u_ppwm/u_ex/_0049_ ),
    .C(\u_ppwm/u_ex/_0050_ ),
    .A(net446),
    .Y(\u_ppwm/u_ex/_0057_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net369));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0607_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net218),
    .A2(\u_ppwm/u_ex/_0057_ ),
    .Y(\u_ppwm/u_ex/_0001_ ),
    .B1(\u_ppwm/u_ex/_0032_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0608_  (.Y(\u_ppwm/u_ex/_0058_ ),
    .B(\u_ppwm/instr[1] ),
    .A_N(\u_ppwm/u_ex/cmp_flag_q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 \u_ppwm/u_ex/_0609_  (.X(\u_ppwm/u_ex/_0059_ ),
    .A(net388),
    .B(\u_ppwm/instr[0] ),
    .C(\u_ppwm/u_ex/_0058_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_ex/_0610_  (.B(\u_ppwm/instr[0] ),
    .C(\u_ppwm/u_ex/_0058_ ),
    .A(\u_ppwm/instr[2] ),
    .Y(\u_ppwm/u_ex/_0060_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0611_  (.B1(net446),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0061_ ),
    .VSS(VGND),
    .A1(net385),
    .A2(\u_ppwm/u_ex/_0060_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0612_  (.B(\u_ppwm/u_ex/_0061_ ),
    .A(net483),
    .X(\u_ppwm/u_ex/_0062_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0613_  (.A(\u_ppwm/u_ex/_0032_ ),
    .B(\u_ppwm/u_ex/_0062_ ),
    .Y(\u_ppwm/u_ex/_0003_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0614_  (.B1(net447),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0063_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0046_ ),
    .A2(\u_ppwm/u_ex/_0059_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0615_  (.B1(\u_ppwm/u_ex/_0063_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0064_ ),
    .VSS(VGND),
    .A1(net473),
    .A2(net483));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0616_  (.B(net383),
    .A(net473),
    .X(\u_ppwm/u_ex/_0065_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0617_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net483),
    .A2(net385),
    .Y(\u_ppwm/u_ex/_0066_ ),
    .B1(\u_ppwm/u_ex/_0065_ ));
 sg13g2_and3_1 \u_ppwm/u_ex/_0618_  (.X(\u_ppwm/u_ex/_0067_ ),
    .A(net483),
    .B(net385),
    .C(\u_ppwm/u_ex/_0065_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 \u_ppwm/u_ex/_0619_  (.A(\u_ppwm/u_ex/_0060_ ),
    .B(\u_ppwm/u_ex/_0066_ ),
    .C(\u_ppwm/u_ex/_0067_ ),
    .X(\u_ppwm/u_ex/_0068_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0620_  (.B1(net512),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0069_ ),
    .VSS(VGND),
    .A1(net447),
    .A2(net473));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0621_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0064_ ),
    .A2(\u_ppwm/u_ex/_0068_ ),
    .Y(\u_ppwm/u_ex/_0004_ ),
    .B1(\u_ppwm/u_ex/_0069_ ));
 sg13g2_or2_1 \u_ppwm/u_ex/_0622_  (.VSS(VGND),
    .VDD(VPWR),
    .X(\u_ppwm/u_ex/_0070_ ),
    .B(\u_ppwm/u_ex/_0046_ ),
    .A(net469));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0623_  (.A(net469),
    .B(\u_ppwm/u_ex/_0059_ ),
    .Y(\u_ppwm/u_ex/_0071_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0624_  (.B1(\u_ppwm/u_ex/_0070_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0072_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0063_ ),
    .A2(\u_ppwm/u_ex/_0071_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0625_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net473),
    .A2(net383),
    .Y(\u_ppwm/u_ex/_0073_ ),
    .B1(\u_ppwm/u_ex/_0067_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0626_  (.Y(\u_ppwm/u_ex/_0074_ ),
    .A(net469),
    .B(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0627_  (.Y(\u_ppwm/u_ex/_0075_ ),
    .A(net469),
    .B(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0628_  (.Y(\u_ppwm/u_ex/_0076_ ),
    .A(\u_ppwm/u_ex/_0073_ ),
    .B(\u_ppwm/u_ex/_0075_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0629_  (.B1(\u_ppwm/u_ex/_0072_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0077_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0060_ ),
    .A2(\u_ppwm/u_ex/_0076_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0630_  (.B1(\u_ppwm/u_ex/_0077_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0078_ ),
    .VSS(VGND),
    .A1(net447),
    .A2(net469));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0631_  (.A(\u_ppwm/u_ex/_0032_ ),
    .B(net674),
    .Y(\u_ppwm/u_ex/_0005_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0632_  (.B1(\u_ppwm/u_ex/_0074_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0079_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0073_ ),
    .A2(\u_ppwm/u_ex/_0075_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0633_  (.Y(\u_ppwm/u_ex/_0080_ ),
    .A(net468),
    .B(net375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0634_  (.Y(\u_ppwm/u_ex/_0081_ ),
    .A(\u_ppwm/u_ex/_0079_ ),
    .B(\u_ppwm/u_ex/_0080_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0635_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net469),
    .A2(\u_ppwm/u_ex/_0046_ ),
    .Y(\u_ppwm/u_ex/_0082_ ),
    .B1(net468));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0636_  (.Y(\u_ppwm/u_ex/_0083_ ),
    .A(\u_ppwm/u_ex/_0047_ ),
    .B(\u_ppwm/u_ex/_0060_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0637_  (.B1(net447),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0084_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0082_ ),
    .A2(\u_ppwm/u_ex/_0083_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0638_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0059_ ),
    .A2(\u_ppwm/u_ex/_0081_ ),
    .Y(\u_ppwm/u_ex/_0085_ ),
    .B1(\u_ppwm/u_ex/_0084_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0639_  (.B1(net501),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0086_ ),
    .VSS(VGND),
    .A1(net468),
    .A2(net447));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0640_  (.A(\u_ppwm/u_ex/_0085_ ),
    .B(net684),
    .Y(\u_ppwm/u_ex/_0006_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0641_  (.Y(\u_ppwm/u_ex/_0087_ ),
    .A(\u_ppwm/u_ex/_0524_ ),
    .B(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0642_  (.Y(\u_ppwm/u_ex/_0088_ ),
    .B1(\u_ppwm/global_counter[4] ),
    .B2(\u_ppwm/u_ex/_0528_ ),
    .A2(\u_ppwm/global_counter[5] ),
    .A1(\u_ppwm/u_ex/_0527_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0643_  (.Y(\u_ppwm/u_ex/_0089_ ),
    .B(net444),
    .A_N(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0644_  (.A(net445),
    .B_N(\u_ppwm/u_ex/reg_value_q[0] ),
    .Y(\u_ppwm/u_ex/_0090_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0645_  (.A(net444),
    .B_N(net453),
    .Y(\u_ppwm/u_ex/_0091_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0646_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0090_ ),
    .C1(\u_ppwm/u_ex/_0091_ ),
    .B1(\u_ppwm/u_ex/_0089_ ),
    .A1(net451),
    .Y(\u_ppwm/u_ex/_0092_ ),
    .A2(\u_ppwm/u_ex/_0044_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0647_  (.Y(\u_ppwm/u_ex/_0093_ ),
    .B(\u_ppwm/global_counter[3] ),
    .A_N(net450),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0648_  (.B1(\u_ppwm/u_ex/_0093_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0094_ ),
    .VSS(VGND),
    .A1(net452),
    .A2(\u_ppwm/u_ex/_0044_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0649_  (.Y(\u_ppwm/u_ex/_0095_ ),
    .B1(\u_ppwm/u_ex/_0043_ ),
    .B2(net450),
    .A2(\u_ppwm/u_ex/_0042_ ),
    .A1(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0650_  (.B1(\u_ppwm/u_ex/_0095_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0096_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0092_ ),
    .A2(\u_ppwm/u_ex/_0094_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0651_  (.A(\u_ppwm/u_ex/_0527_ ),
    .B(\u_ppwm/global_counter[5] ),
    .Y(\u_ppwm/u_ex/_0097_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0652_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0096_ ),
    .C1(\u_ppwm/u_ex/_0097_ ),
    .B1(\u_ppwm/u_ex/_0088_ ),
    .A1(net448),
    .Y(\u_ppwm/u_ex/_0098_ ),
    .A2(\u_ppwm/u_ex/_0041_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0653_  (.Y(\u_ppwm/u_ex/_0099_ ),
    .A(\u_ppwm/u_ex/_0525_ ),
    .B(\u_ppwm/global_counter[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0654_  (.B1(\u_ppwm/u_ex/_0099_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0100_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/reg_value_q[6] ),
    .A2(\u_ppwm/u_ex/_0041_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0655_  (.Y(\u_ppwm/u_ex/_0101_ ),
    .B(\u_ppwm/u_ex/reg_value_q[8] ),
    .A_N(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0656_  (.B1(\u_ppwm/u_ex/_0101_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0102_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0525_ ),
    .A2(\u_ppwm/global_counter[7] ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0657_  (.B(net441),
    .A(\u_ppwm/u_ex/reg_value_q[9] ),
    .X(\u_ppwm/u_ex/_0103_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0658_  (.A(\u_ppwm/u_ex/_0087_ ),
    .B(\u_ppwm/u_ex/_0103_ ),
    .Y(\u_ppwm/u_ex/_0104_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0659_  (.Y(\u_ppwm/u_ex/_0105_ ),
    .B(\u_ppwm/u_ex/_0087_ ),
    .A_N(\u_ppwm/u_ex/_0102_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0660_  (.A(\u_ppwm/u_ex/_0103_ ),
    .B(\u_ppwm/u_ex/_0105_ ),
    .Y(\u_ppwm/u_ex/_0106_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0661_  (.B1(\u_ppwm/u_ex/_0106_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0107_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0098_ ),
    .A2(\u_ppwm/u_ex/_0100_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0662_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0523_ ),
    .A2(net441),
    .Y(\u_ppwm/u_ex/_0108_ ),
    .B1(\u_ppwm/u_ex/_0104_ ));
 sg13g2_and4_1 \u_ppwm/u_ex/_0663_  (.A(net370),
    .B(\u_ppwm/u_ex/_0050_ ),
    .C(\u_ppwm/u_ex/_0107_ ),
    .D(\u_ppwm/u_ex/_0108_ ),
    .X(\u_ppwm/u_ex/_0109_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0664_  (.A(net439),
    .B_N(net456),
    .Y(\u_ppwm/u_ex/_0110_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0665_  (.A(net464),
    .B_N(\u_ppwm/global_counter[11] ),
    .Y(\u_ppwm/u_ex/_0111_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0666_  (.Y(\u_ppwm/u_ex/_0112_ ),
    .B(net466),
    .A_N(\u_ppwm/global_counter[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0667_  (.Y(\u_ppwm/u_ex/_0113_ ),
    .B(net462),
    .A_N(\u_ppwm/global_counter[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0668_  (.B1(\u_ppwm/u_ex/_0113_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0114_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0030_ ),
    .A2(net440));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0669_  (.Y(\u_ppwm/u_ex/_0115_ ),
    .B(net464),
    .A_N(\u_ppwm/global_counter[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0670_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0112_ ),
    .A2(\u_ppwm/u_ex/_0115_ ),
    .Y(\u_ppwm/u_ex/_0116_ ),
    .B1(\u_ppwm/u_ex/_0111_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0671_  (.Y(\u_ppwm/u_ex/_0117_ ),
    .B1(net440),
    .B2(\u_ppwm/u_ex/_0030_ ),
    .A2(\u_ppwm/global_counter[13] ),
    .A1(\u_ppwm/u_ex/_0029_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0672_  (.B1(\u_ppwm/u_ex/_0117_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0118_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0114_ ),
    .A2(\u_ppwm/u_ex/_0116_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0673_  (.A(net463),
    .B(\u_ppwm/u_ex/_0040_ ),
    .C(\u_ppwm/u_ex/_0113_ ),
    .Y(\u_ppwm/u_ex/_0119_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0674_  (.Y(\u_ppwm/u_ex/_0120_ ),
    .B(\u_ppwm/global_counter[15] ),
    .A_N(net458),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0675_  (.B1(\u_ppwm/u_ex/_0120_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0121_ ),
    .VSS(VGND),
    .A1(net460),
    .A2(\u_ppwm/u_ex/_0039_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0676_  (.Y(\u_ppwm/u_ex/_0122_ ),
    .B(net458),
    .A_N(\u_ppwm/global_counter[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0677_  (.B1(\u_ppwm/u_ex/_0122_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0123_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0534_ ),
    .A2(\u_ppwm/global_counter[14] ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0678_  (.A(\u_ppwm/u_ex/_0119_ ),
    .B(\u_ppwm/u_ex/_0121_ ),
    .C(\u_ppwm/u_ex/_0123_ ),
    .Y(\u_ppwm/u_ex/_0124_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0679_  (.A(net457),
    .B_N(net439),
    .Y(\u_ppwm/u_ex/_0125_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0680_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0118_ ),
    .C1(\u_ppwm/u_ex/_0125_ ),
    .B1(\u_ppwm/u_ex/_0124_ ),
    .A1(\u_ppwm/u_ex/_0121_ ),
    .Y(\u_ppwm/u_ex/_0126_ ),
    .A2(\u_ppwm/u_ex/_0122_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0681_  (.Y(\u_ppwm/u_ex/_0127_ ),
    .A(\u_ppwm/u_ex/_0532_ ),
    .B(\u_ppwm/global_counter[17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0682_  (.B1(\u_ppwm/u_ex/_0127_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0128_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0110_ ),
    .A2(\u_ppwm/u_ex/_0126_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0683_  (.Y(\u_ppwm/u_ex/_0129_ ),
    .A(\u_ppwm/u_ex/_0530_ ),
    .B(\u_ppwm/global_counter[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0684_  (.B1(\u_ppwm/u_ex/_0129_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0130_ ),
    .VSS(VGND),
    .A1(net455),
    .A2(\u_ppwm/u_ex/_0038_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0685_  (.A(\u_ppwm/u_ex/_0531_ ),
    .B(\u_ppwm/global_counter[18] ),
    .Y(\u_ppwm/u_ex/_0131_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0686_  (.Y(\u_ppwm/u_ex/_0132_ ),
    .B(net454),
    .A_N(\u_ppwm/global_counter[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0687_  (.B1(\u_ppwm/u_ex/_0132_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0133_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0532_ ),
    .A2(\u_ppwm/global_counter[17] ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0688_  (.A(\u_ppwm/u_ex/_0130_ ),
    .B(\u_ppwm/u_ex/_0131_ ),
    .C(\u_ppwm/u_ex/_0133_ ),
    .Y(\u_ppwm/u_ex/_0134_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0689_  (.A(net381),
    .B(net385),
    .Y(\u_ppwm/u_ex/_0135_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_ex/_0690_  (.A(net379),
    .B(\u_ppwm/u_ex/_0135_ ),
    .X(\u_ppwm/u_ex/_0136_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0691_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0137_ ),
    .A(net366),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0692_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0128_ ),
    .C1(\u_ppwm/u_ex/_0137_ ),
    .B1(\u_ppwm/u_ex/_0134_ ),
    .A1(\u_ppwm/u_ex/_0130_ ),
    .Y(\u_ppwm/u_ex/_0138_ ),
    .A2(\u_ppwm/u_ex/_0132_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0693_  (.Y(\u_ppwm/u_ex/_0139_ ),
    .A(\u_ppwm/u_ex/reg_value_q[4] ),
    .B(\u_ppwm/u_ex/_0039_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0694_  (.A(\u_ppwm/u_ex/reg_value_q[1] ),
    .B_N(\u_ppwm/global_counter[11] ),
    .Y(\u_ppwm/u_ex/_0140_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0695_  (.Y(\u_ppwm/u_ex/_0141_ ),
    .B(\u_ppwm/u_ex/reg_value_q[0] ),
    .A_N(\u_ppwm/global_counter[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0696_  (.Y(\u_ppwm/u_ex/_0142_ ),
    .B(net450),
    .A_N(\u_ppwm/global_counter[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0697_  (.B1(\u_ppwm/u_ex/_0142_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0143_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0529_ ),
    .A2(net440));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0698_  (.Y(\u_ppwm/u_ex/_0144_ ),
    .B(\u_ppwm/u_ex/reg_value_q[1] ),
    .A_N(\u_ppwm/global_counter[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0699_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0141_ ),
    .A2(\u_ppwm/u_ex/_0144_ ),
    .Y(\u_ppwm/u_ex/_0145_ ),
    .B1(\u_ppwm/u_ex/_0140_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0700_  (.A(net452),
    .B_N(net440),
    .Y(\u_ppwm/u_ex/_0146_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0701_  (.A(\u_ppwm/u_ex/reg_value_q[3] ),
    .B_N(\u_ppwm/global_counter[13] ),
    .Y(\u_ppwm/u_ex/_0147_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0702_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0146_ ),
    .C1(\u_ppwm/u_ex/_0147_ ),
    .B1(\u_ppwm/u_ex/_0142_ ),
    .A1(\u_ppwm/u_ex/_0528_ ),
    .Y(\u_ppwm/u_ex/_0148_ ),
    .A2(\u_ppwm/global_counter[14] ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0703_  (.B1(\u_ppwm/u_ex/_0148_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0149_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0143_ ),
    .A2(\u_ppwm/u_ex/_0145_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0704_  (.Y(\u_ppwm/u_ex/_0150_ ),
    .B1(\u_ppwm/u_ex/_0139_ ),
    .B2(\u_ppwm/u_ex/_0149_ ),
    .A2(\u_ppwm/global_counter[15] ),
    .A1(\u_ppwm/u_ex/_0527_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0705_  (.Y(\u_ppwm/u_ex/_0151_ ),
    .B(net448),
    .A_N(net439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0706_  (.B1(\u_ppwm/u_ex/_0151_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0152_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0527_ ),
    .A2(\u_ppwm/global_counter[15] ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0707_  (.Y(\u_ppwm/u_ex/_0153_ ),
    .B1(net439),
    .B2(\u_ppwm/u_ex/_0526_ ),
    .A2(\u_ppwm/global_counter[17] ),
    .A1(\u_ppwm/u_ex/_0525_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0708_  (.B1(\u_ppwm/u_ex/_0153_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0154_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0150_ ),
    .A2(\u_ppwm/u_ex/_0152_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0709_  (.Y(\u_ppwm/u_ex/_0155_ ),
    .A(\u_ppwm/u_ex/_0523_ ),
    .B(\u_ppwm/global_counter[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0710_  (.B1(\u_ppwm/u_ex/_0155_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0156_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/reg_value_q[8] ),
    .A2(\u_ppwm/u_ex/_0038_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0711_  (.A(\u_ppwm/u_ex/_0524_ ),
    .B(\u_ppwm/global_counter[18] ),
    .Y(\u_ppwm/u_ex/_0157_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0712_  (.Y(\u_ppwm/u_ex/_0158_ ),
    .B(\u_ppwm/u_ex/reg_value_q[9] ),
    .A_N(\u_ppwm/global_counter[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0713_  (.B1(\u_ppwm/u_ex/_0158_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0159_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0525_ ),
    .A2(\u_ppwm/global_counter[17] ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0714_  (.A(\u_ppwm/u_ex/_0156_ ),
    .B(\u_ppwm/u_ex/_0157_ ),
    .C(\u_ppwm/u_ex/_0159_ ),
    .Y(\u_ppwm/u_ex/_0160_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_ex/_0715_  (.A(net377),
    .B(\u_ppwm/u_ex/_0050_ ),
    .X(\u_ppwm/u_ex/_0161_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0716_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0162_ ),
    .A(net364),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0717_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0154_ ),
    .C1(\u_ppwm/u_ex/_0162_ ),
    .B1(\u_ppwm/u_ex/_0160_ ),
    .A1(\u_ppwm/u_ex/_0156_ ),
    .Y(\u_ppwm/u_ex/_0163_ ),
    .A2(\u_ppwm/u_ex/_0158_ ));
 sg13g2_and4_1 \u_ppwm/u_ex/_0718_  (.A(net446),
    .B(net388),
    .C(\u_ppwm/u_ex/_0033_ ),
    .D(\u_ppwm/instr[1] ),
    .X(\u_ppwm/u_ex/_0164_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0719_  (.A(\u_ppwm/u_ex/_0526_ ),
    .B(net457),
    .Y(\u_ppwm/u_ex/_0165_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0720_  (.Y(\u_ppwm/u_ex/_0166_ ),
    .B(net465),
    .A_N(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0721_  (.A(net466),
    .B_N(\u_ppwm/u_ex/reg_value_q[0] ),
    .Y(\u_ppwm/u_ex/_0167_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0722_  (.A(net465),
    .B_N(net453),
    .Y(\u_ppwm/u_ex/_0168_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0723_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0167_ ),
    .C1(\u_ppwm/u_ex/_0168_ ),
    .B1(\u_ppwm/u_ex/_0166_ ),
    .A1(net452),
    .Y(\u_ppwm/u_ex/_0169_ ),
    .A2(\u_ppwm/u_ex/_0030_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0724_  (.Y(\u_ppwm/u_ex/_0170_ ),
    .B(net462),
    .A_N(\u_ppwm/u_ex/reg_value_q[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0725_  (.B1(\u_ppwm/u_ex/_0170_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0171_ ),
    .VSS(VGND),
    .A1(net452),
    .A2(\u_ppwm/u_ex/_0030_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0726_  (.A(\u_ppwm/u_ex/reg_value_q[5] ),
    .B_N(net459),
    .Y(\u_ppwm/u_ex/_0172_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0727_  (.A(net459),
    .B_N(\u_ppwm/u_ex/reg_value_q[5] ),
    .Y(\u_ppwm/u_ex/_0173_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0728_  (.A(net462),
    .B_N(\u_ppwm/u_ex/reg_value_q[3] ),
    .Y(\u_ppwm/u_ex/_0174_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0729_  (.B(net460),
    .A(net449),
    .X(\u_ppwm/u_ex/_0175_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 \u_ppwm/u_ex/_0730_  (.A(\u_ppwm/u_ex/_0172_ ),
    .B(\u_ppwm/u_ex/_0173_ ),
    .C(\u_ppwm/u_ex/_0174_ ),
    .D(\u_ppwm/u_ex/_0175_ ),
    .Y(\u_ppwm/u_ex/_0176_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0731_  (.B1(\u_ppwm/u_ex/_0176_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0177_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0169_ ),
    .A2(\u_ppwm/u_ex/_0171_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0732_  (.A(net449),
    .B(\u_ppwm/u_ex/_0534_ ),
    .C(\u_ppwm/u_ex/_0173_ ),
    .Y(\u_ppwm/u_ex/_0178_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0733_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0527_ ),
    .C1(\u_ppwm/u_ex/_0178_ ),
    .B1(net458),
    .A1(\u_ppwm/u_ex/_0526_ ),
    .Y(\u_ppwm/u_ex/_0179_ ),
    .A2(net457));
 sg13g2_a21o_1 \u_ppwm/u_ex/_0734_  (.A2(\u_ppwm/u_ex/_0179_ ),
    .A1(\u_ppwm/u_ex/_0177_ ),
    .B1(\u_ppwm/u_ex/_0165_ ),
    .X(\u_ppwm/u_ex/_0180_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0735_  (.Y(\u_ppwm/u_ex/_0181_ ),
    .A(\u_ppwm/u_ex/_0525_ ),
    .B(\u_ppwm/pwm_value[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0736_  (.Y(\u_ppwm/u_ex/_0182_ ),
    .B1(net455),
    .B2(\u_ppwm/u_ex/_0524_ ),
    .A2(net454),
    .A1(\u_ppwm/u_ex/_0523_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0737_  (.A(\u_ppwm/u_ex/_0523_ ),
    .B(net454),
    .Y(\u_ppwm/u_ex/_0183_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0738_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/reg_value_q[7] ),
    .C1(\u_ppwm/u_ex/_0183_ ),
    .B1(\u_ppwm/u_ex/_0532_ ),
    .A1(\u_ppwm/u_ex/reg_value_q[8] ),
    .Y(\u_ppwm/u_ex/_0184_ ),
    .A2(\u_ppwm/u_ex/_0531_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0739_  (.Y(\u_ppwm/u_ex/_0185_ ),
    .A(\u_ppwm/u_ex/_0182_ ),
    .B(\u_ppwm/u_ex/_0184_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0740_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0180_ ),
    .A2(\u_ppwm/u_ex/_0181_ ),
    .Y(\u_ppwm/u_ex/_0186_ ),
    .B1(\u_ppwm/u_ex/_0185_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0741_  (.Y(\u_ppwm/u_ex/_0187_ ),
    .A(net382),
    .B(net370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 \u_ppwm/u_ex/_0742_  (.A(net387),
    .B(net363),
    .Y(\u_ppwm/u_ex/_0188_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0743_  (.B1(net356),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0189_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0182_ ),
    .A2(\u_ppwm/u_ex/_0183_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0744_  (.B1(\u_ppwm/u_ex/_0164_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0190_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0186_ ),
    .A2(\u_ppwm/u_ex/_0189_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0745_  (.A(net464),
    .B_N(net444),
    .Y(\u_ppwm/u_ex/_0191_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0746_  (.Y(\u_ppwm/u_ex/_0192_ ),
    .B(net466),
    .A_N(net445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0747_  (.Y(\u_ppwm/u_ex/_0193_ ),
    .B(net462),
    .A_N(\u_ppwm/global_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0748_  (.B1(\u_ppwm/u_ex/_0193_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0194_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0030_ ),
    .A2(net443));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0749_  (.Y(\u_ppwm/u_ex/_0195_ ),
    .B(net464),
    .A_N(net444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0750_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0192_ ),
    .A2(\u_ppwm/u_ex/_0195_ ),
    .Y(\u_ppwm/u_ex/_0196_ ),
    .B1(\u_ppwm/u_ex/_0191_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0751_  (.Y(\u_ppwm/u_ex/_0197_ ),
    .B1(net443),
    .B2(\u_ppwm/u_ex/_0030_ ),
    .A2(\u_ppwm/global_counter[3] ),
    .A1(\u_ppwm/u_ex/_0029_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0752_  (.B1(\u_ppwm/u_ex/_0197_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0198_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0194_ ),
    .A2(\u_ppwm/u_ex/_0196_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0753_  (.A(net463),
    .B(\u_ppwm/u_ex/_0193_ ),
    .Y(\u_ppwm/u_ex/_0199_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0754_  (.Y(\u_ppwm/u_ex/_0200_ ),
    .B1(net443),
    .B2(\u_ppwm/u_ex/_0199_ ),
    .A2(\u_ppwm/u_ex/_0042_ ),
    .A1(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0755_  (.A(net461),
    .B(\u_ppwm/u_ex/_0042_ ),
    .Y(\u_ppwm/u_ex/_0201_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0756_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0200_ ),
    .C1(\u_ppwm/u_ex/_0201_ ),
    .B1(\u_ppwm/u_ex/_0198_ ),
    .A1(\u_ppwm/u_ex/_0533_ ),
    .Y(\u_ppwm/u_ex/_0202_ ),
    .A2(\u_ppwm/global_counter[5] ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0757_  (.A(\u_ppwm/u_ex/_0532_ ),
    .B(\u_ppwm/global_counter[7] ),
    .Y(\u_ppwm/u_ex/_0203_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0758_  (.A(\u_ppwm/u_ex/_0533_ ),
    .B(\u_ppwm/global_counter[5] ),
    .Y(\u_ppwm/u_ex/_0204_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0759_  (.B(\u_ppwm/global_counter[6] ),
    .A(net456),
    .X(\u_ppwm/u_ex/_0205_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 \u_ppwm/u_ex/_0760_  (.A(\u_ppwm/u_ex/_0202_ ),
    .B(\u_ppwm/u_ex/_0203_ ),
    .C(\u_ppwm/u_ex/_0204_ ),
    .D(\u_ppwm/u_ex/_0205_ ),
    .Y(\u_ppwm/u_ex/_0206_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0761_  (.A(net457),
    .B(\u_ppwm/u_ex/_0041_ ),
    .C(\u_ppwm/u_ex/_0203_ ),
    .Y(\u_ppwm/u_ex/_0207_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0762_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0532_ ),
    .C1(\u_ppwm/u_ex/_0207_ ),
    .B1(\u_ppwm/global_counter[7] ),
    .A1(\u_ppwm/u_ex/_0531_ ),
    .Y(\u_ppwm/u_ex/_0208_ ),
    .A2(net442));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0763_  (.A(\u_ppwm/u_ex/_0206_ ),
    .B_N(\u_ppwm/u_ex/_0208_ ),
    .Y(\u_ppwm/u_ex/_0209_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0764_  (.Y(\u_ppwm/u_ex/_0210_ ),
    .B(net455),
    .A_N(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0765_  (.B1(\u_ppwm/u_ex/_0210_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0211_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0530_ ),
    .A2(net441));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0766_  (.A(net454),
    .B_N(net441),
    .Y(\u_ppwm/u_ex/_0212_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 \u_ppwm/u_ex/_0767_  (.A(net382),
    .B(net386),
    .C(net378),
    .D(\u_ppwm/u_ex/_0212_ ),
    .Y(\u_ppwm/u_ex/_0213_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0768_  (.B1(\u_ppwm/u_ex/_0213_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0214_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0209_ ),
    .A2(\u_ppwm/u_ex/_0211_ ));
 sg13g2_nor4_1 \u_ppwm/u_ex/_0769_  (.A(\u_ppwm/u_ex/_0109_ ),
    .B(\u_ppwm/u_ex/_0138_ ),
    .C(\u_ppwm/u_ex/_0163_ ),
    .D(\u_ppwm/u_ex/_0190_ ),
    .Y(\u_ppwm/u_ex/_0215_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0770_  (.B1(net492),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0216_ ),
    .VSS(VGND),
    .A1(net648),
    .A2(\u_ppwm/u_ex/_0164_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0771_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0214_ ),
    .A2(\u_ppwm/u_ex/_0215_ ),
    .Y(\u_ppwm/u_ex/_0007_ ),
    .B1(net649));
 sg13g2_nand4_1 \u_ppwm/u_ex/_0772_  (.B(net383),
    .C(\u_ppwm/u_ex/_0049_ ),
    .A(net446),
    .Y(\u_ppwm/u_ex/_0217_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net369));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0773_  (.B1(net492),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0218_ ),
    .VSS(VGND),
    .A1(net384),
    .A2(\u_ppwm/u_ex/_0217_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0774_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0031_ ),
    .A2(\u_ppwm/u_ex/_0217_ ),
    .Y(\u_ppwm/u_ex/_0008_ ),
    .B1(\u_ppwm/u_ex/_0218_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_0775_  (.A(net388),
    .B(\u_ppwm/u_ex/_0048_ ),
    .X(\u_ppwm/u_ex/_0219_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \u_ppwm/u_ex/_0776_  (.Y(\u_ppwm/u_ex/_0220_ ),
    .A(net388),
    .B(\u_ppwm/u_ex/_0048_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 \u_ppwm/u_ex/_0777_  (.A(net366),
    .B(net364),
    .C(net359),
    .Y(\u_ppwm/u_ex/_0221_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0778_  (.Y(\u_ppwm/u_ex/_0222_ ),
    .B1(net365),
    .B2(net575),
    .A2(net366),
    .A1(net445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 \u_ppwm/u_ex/_0779_  (.A(net388),
    .B_N(\u_ppwm/instr[1] ),
    .Y(\u_ppwm/u_ex/_0223_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_ex/_0780_  (.A(\u_ppwm/u_ex/_0033_ ),
    .B(\u_ppwm/u_ex/_0223_ ),
    .X(\u_ppwm/u_ex/_0224_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0781_  (.Y(\u_ppwm/u_ex/_0225_ ),
    .A(\u_ppwm/u_ex/_0033_ ),
    .B(\u_ppwm/u_ex/_0223_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0782_  (.Y(\u_ppwm/u_ex/_0226_ ),
    .A(net466),
    .B(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0783_  (.B(net383),
    .A(net466),
    .X(\u_ppwm/u_ex/_0227_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 \u_ppwm/u_ex/_0784_  (.A(\u_ppwm/u_ex/_0219_ ),
    .B(\u_ppwm/u_ex/_0223_ ),
    .Y(\u_ppwm/u_ex/_0228_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0785_  (.Y(\u_ppwm/u_ex/_0229_ ),
    .B1(\u_ppwm/u_ex/_0228_ ),
    .B2(net382),
    .A2(\u_ppwm/u_ex/_0227_ ),
    .A1(\u_ppwm/u_ex/_0224_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0786_  (.B1(\u_ppwm/u_ex/_0229_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0230_ ),
    .VSS(VGND),
    .A1(net359),
    .A2(\u_ppwm/u_ex/_0222_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0787_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net660),
    .A2(\u_ppwm/u_ex/_0221_ ),
    .Y(\u_ppwm/u_ex/_0231_ ),
    .B1(\u_ppwm/u_ex/_0230_ ));
 sg13g2_nand2_2 \u_ppwm/u_ex/_0788_  (.Y(\u_ppwm/u_ex/_0232_ ),
    .A(\u_ppwm/instr[0] ),
    .B(\u_ppwm/u_ex/_0223_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0789_  (.A(net381),
    .B(net375),
    .Y(\u_ppwm/u_ex/_0233_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 \u_ppwm/u_ex/_0790_  (.A(\u_ppwm/u_ex/_0232_ ),
    .B_N(\u_ppwm/u_ex/_0233_ ),
    .Y(\u_ppwm/u_ex/_0234_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 \u_ppwm/u_ex/_0791_  (.VSS(VGND),
    .VDD(VPWR),
    .X(\u_ppwm/u_ex/_0235_ ),
    .B(net386),
    .A(net464));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0792_  (.B1(\u_ppwm/u_ex/_0235_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0236_ ),
    .VSS(VGND),
    .A1(net453),
    .A2(\u_ppwm/u_ex/_0034_ ));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0793_  (.A0(net463),
    .A1(net451),
    .S(net386),
    .X(\u_ppwm/u_ex/_0237_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0794_  (.Y(\u_ppwm/u_ex/_0238_ ),
    .A(net379),
    .B(\u_ppwm/u_ex/_0237_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0795_  (.B1(\u_ppwm/u_ex/_0238_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0239_ ),
    .VSS(VGND),
    .A1(net378),
    .A2(\u_ppwm/u_ex/_0236_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0796_  (.A(net382),
    .B(\u_ppwm/u_ex/_0035_ ),
    .Y(\u_ppwm/u_ex/_0240_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 \u_ppwm/u_ex/_0797_  (.A(\u_ppwm/u_ex/_0232_ ),
    .B_N(\u_ppwm/u_ex/_0240_ ),
    .Y(\u_ppwm/u_ex/_0241_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0798_  (.A0(net461),
    .A1(net449),
    .S(net386),
    .X(\u_ppwm/u_ex/_0242_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0799_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0243_ ),
    .A(\u_ppwm/u_ex/_0242_ ),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0800_  (.A0(net462),
    .A1(net450),
    .S(net386),
    .X(\u_ppwm/u_ex/_0244_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0801_  (.A0(\u_ppwm/u_ex/_0242_ ),
    .A1(\u_ppwm/u_ex/_0244_ ),
    .S(net370),
    .X(\u_ppwm/u_ex/_0245_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0802_  (.Y(\u_ppwm/u_ex/_0246_ ),
    .B1(\u_ppwm/u_ex/_0241_ ),
    .B2(\u_ppwm/u_ex/_0245_ ),
    .A2(\u_ppwm/u_ex/_0239_ ),
    .A1(\u_ppwm/u_ex/_0234_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 \u_ppwm/u_ex/_0803_  (.A(\u_ppwm/u_ex/_0135_ ),
    .B(net364),
    .C(net361),
    .X(\u_ppwm/u_ex/_0247_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0804_  (.A(net388),
    .B(\u_ppwm/u_ex/_0048_ ),
    .Y(\u_ppwm/u_ex/_0248_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0805_  (.A(net388),
    .B(net385),
    .C(\u_ppwm/u_ex/_0048_ ),
    .Y(\u_ppwm/u_ex/_0249_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0806_  (.B1(net446),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0250_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0219_ ),
    .A2(\u_ppwm/u_ex/_0249_ ));
 sg13g2_nor2b_2 \u_ppwm/u_ex/_0807_  (.A(\u_ppwm/u_ex/_0250_ ),
    .B_N(\u_ppwm/u_ex/_0247_ ),
    .Y(\u_ppwm/u_ex/_0251_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_ex/_0808_  (.A(\u_ppwm/u_ex/_0246_ ),
    .B(net354),
    .X(\u_ppwm/u_ex/_0252_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0809_  (.B1(net506),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0253_ ),
    .VSS(VGND),
    .A1(net466),
    .A2(net354));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0810_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0231_ ),
    .A2(\u_ppwm/u_ex/_0252_ ),
    .Y(\u_ppwm/u_ex/_0009_ ),
    .B1(\u_ppwm/u_ex/_0253_ ));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0811_  (.A0(net459),
    .A1(\u_ppwm/u_ex/reg_value_q[5] ),
    .S(net386),
    .X(\u_ppwm/u_ex/_0254_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0812_  (.A0(\u_ppwm/u_ex/_0527_ ),
    .A1(\u_ppwm/u_ex/_0533_ ),
    .S(\u_ppwm/u_ex/_0034_ ),
    .X(\u_ppwm/u_ex/_0255_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0813_  (.A0(\u_ppwm/u_ex/_0242_ ),
    .A1(\u_ppwm/u_ex/_0254_ ),
    .S(net377),
    .X(\u_ppwm/u_ex/_0256_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_0814_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0257_ ),
    .A(\u_ppwm/u_ex/_0256_ ),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0815_  (.A0(net466),
    .A1(\u_ppwm/u_ex/reg_value_q[0] ),
    .S(net386),
    .X(\u_ppwm/u_ex/_0258_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0816_  (.Y(\u_ppwm/u_ex/_0259_ ),
    .A(net370),
    .B(\u_ppwm/u_ex/_0258_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0817_  (.B1(\u_ppwm/u_ex/_0259_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0260_ ),
    .VSS(VGND),
    .A1(net370),
    .A2(\u_ppwm/u_ex/_0236_ ));
 sg13g2_and3_2 \u_ppwm/u_ex/_0818_  (.X(\u_ppwm/u_ex/_0261_ ),
    .A(\u_ppwm/instr[0] ),
    .B(net381),
    .C(\u_ppwm/u_ex/_0223_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_ex/_0819_  (.B(net381),
    .C(\u_ppwm/u_ex/_0223_ ),
    .A(\u_ppwm/instr[0] ),
    .Y(\u_ppwm/u_ex/_0262_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_ex/_0820_  (.B(\u_ppwm/u_ex/_0260_ ),
    .C(\u_ppwm/u_ex/_0261_ ),
    .A(net369),
    .Y(\u_ppwm/u_ex/_0263_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0821_  (.A0(\u_ppwm/u_ex/_0237_ ),
    .A1(\u_ppwm/u_ex/_0244_ ),
    .S(net378),
    .X(\u_ppwm/u_ex/_0264_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0822_  (.Y(\u_ppwm/u_ex/_0265_ ),
    .B1(\u_ppwm/u_ex/_0264_ ),
    .B2(\u_ppwm/u_ex/_0234_ ),
    .A2(\u_ppwm/u_ex/_0256_ ),
    .A1(\u_ppwm/u_ex/_0241_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0823_  (.Y(\u_ppwm/u_ex/_0266_ ),
    .A(\u_ppwm/u_ex/_0263_ ),
    .B(\u_ppwm/u_ex/_0265_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0824_  (.Y(\u_ppwm/u_ex/_0267_ ),
    .A(net379),
    .B(\u_ppwm/u_ex/_0228_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0825_  (.Y(\u_ppwm/u_ex/_0268_ ),
    .A(net464),
    .B(net379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0826_  (.Y(\u_ppwm/u_ex/_0269_ ),
    .A(net464),
    .B(net379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0827_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0226_ ),
    .A2(\u_ppwm/u_ex/_0269_ ),
    .Y(\u_ppwm/u_ex/_0270_ ),
    .B1(net358));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0828_  (.B1(\u_ppwm/u_ex/_0270_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0271_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0226_ ),
    .A2(\u_ppwm/u_ex/_0269_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_0829_  (.B(\u_ppwm/u_ex/_0267_ ),
    .C(\u_ppwm/u_ex/_0271_ ),
    .A(net354),
    .Y(\u_ppwm/u_ex/_0272_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0830_  (.Y(\u_ppwm/u_ex/_0273_ ),
    .B1(net365),
    .B2(\u_ppwm/global_counter[11] ),
    .A2(net366),
    .A1(net444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0831_  (.Y(\u_ppwm/u_ex/_0274_ ),
    .A(net678),
    .B(\u_ppwm/u_ex/_0221_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0832_  (.B1(\u_ppwm/u_ex/_0274_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0275_ ),
    .VSS(VGND),
    .A1(net360),
    .A2(\u_ppwm/u_ex/_0273_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0833_  (.A(\u_ppwm/u_ex/_0266_ ),
    .B(\u_ppwm/u_ex/_0272_ ),
    .C(\u_ppwm/u_ex/_0275_ ),
    .Y(\u_ppwm/u_ex/_0276_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0834_  (.B1(net508),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0277_ ),
    .VSS(VGND),
    .A1(net464),
    .A2(net354));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0835_  (.A(\u_ppwm/u_ex/_0276_ ),
    .B(\u_ppwm/u_ex/_0277_ ),
    .Y(\u_ppwm/u_ex/_0010_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_ex/_0836_  (.A(net375),
    .B(net377),
    .X(\u_ppwm/u_ex/_0278_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \u_ppwm/u_ex/_0837_  (.Y(\u_ppwm/u_ex/_0279_ ),
    .A(net375),
    .B(net377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0838_  (.A(net368),
    .B(\u_ppwm/u_ex/_0278_ ),
    .Y(\u_ppwm/u_ex/_0280_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 \u_ppwm/u_ex/_0839_  (.Y(\u_ppwm/u_ex/_0281_ ),
    .B(\u_ppwm/u_ex/_0279_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net368));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0840_  (.A(net375),
    .B(\u_ppwm/u_ex/_0036_ ),
    .Y(\u_ppwm/u_ex/_0282_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0841_  (.Y(\u_ppwm/u_ex/_0283_ ),
    .B1(\u_ppwm/u_ex/_0282_ ),
    .B2(\u_ppwm/u_ex/_0258_ ),
    .A2(\u_ppwm/u_ex/_0281_ ),
    .A1(\u_ppwm/u_ex/_0239_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0842_  (.Y(\u_ppwm/u_ex/_0284_ ),
    .A(net381),
    .B(\u_ppwm/u_ex/_0279_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0843_  (.A(\u_ppwm/u_ex/_0232_ ),
    .B(\u_ppwm/u_ex/_0283_ ),
    .C(\u_ppwm/u_ex/_0284_ ),
    .Y(\u_ppwm/u_ex/_0285_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0844_  (.A0(net456),
    .A1(net448),
    .S(net384),
    .X(\u_ppwm/u_ex/_0286_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0845_  (.Y(\u_ppwm/u_ex/_0287_ ),
    .A(net378),
    .B(\u_ppwm/u_ex/_0286_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0846_  (.B1(\u_ppwm/u_ex/_0287_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0288_ ),
    .VSS(VGND),
    .A1(net378),
    .A2(\u_ppwm/u_ex/_0255_ ));
 sg13g2_inv_1 \u_ppwm/u_ex/_0847_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0289_ ),
    .A(\u_ppwm/u_ex/_0288_ ),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0848_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0241_ ),
    .C1(\u_ppwm/u_ex/_0285_ ),
    .B1(\u_ppwm/u_ex/_0288_ ),
    .A1(\u_ppwm/u_ex/_0234_ ),
    .Y(\u_ppwm/u_ex/_0290_ ),
    .A2(\u_ppwm/u_ex/_0245_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0849_  (.B1(\u_ppwm/u_ex/_0268_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0291_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0226_ ),
    .A2(\u_ppwm/u_ex/_0269_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0850_  (.A(\u_ppwm/u_ex/_0030_ ),
    .B(\u_ppwm/u_ex/_0035_ ),
    .Y(\u_ppwm/u_ex/_0292_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0851_  (.B(net373),
    .A(net463),
    .X(\u_ppwm/u_ex/_0293_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0852_  (.Y(\u_ppwm/u_ex/_0294_ ),
    .A(net463),
    .B(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0853_  (.B1(\u_ppwm/u_ex/_0224_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0295_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0291_ ),
    .A2(\u_ppwm/u_ex/_0293_ ));
 sg13g2_a21o_1 \u_ppwm/u_ex/_0854_  (.A2(\u_ppwm/u_ex/_0293_ ),
    .A1(\u_ppwm/u_ex/_0291_ ),
    .B1(\u_ppwm/u_ex/_0295_ ),
    .X(\u_ppwm/u_ex/_0296_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0855_  (.Y(\u_ppwm/u_ex/_0297_ ),
    .B1(net364),
    .B2(net440),
    .A2(net367),
    .A1(net443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0856_  (.Y(\u_ppwm/u_ex/_0298_ ),
    .A(net375),
    .B(\u_ppwm/u_ex/_0228_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0857_  (.B1(\u_ppwm/u_ex/_0298_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0299_ ),
    .VSS(VGND),
    .A1(net359),
    .A2(\u_ppwm/u_ex/_0297_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0858_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net451),
    .A2(\u_ppwm/u_ex/_0221_ ),
    .Y(\u_ppwm/u_ex/_0300_ ),
    .B1(\u_ppwm/u_ex/_0299_ ));
 sg13g2_nand4_1 \u_ppwm/u_ex/_0859_  (.B(\u_ppwm/u_ex/_0290_ ),
    .C(\u_ppwm/u_ex/_0296_ ),
    .A(net354),
    .Y(\u_ppwm/u_ex/_0301_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0300_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0860_  (.B1(net508),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0302_ ),
    .VSS(VGND),
    .A1(net463),
    .A2(net354));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0861_  (.A(\u_ppwm/u_ex/_0302_ ),
    .B_N(\u_ppwm/u_ex/_0301_ ),
    .Y(\u_ppwm/u_ex/_0011_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0862_  (.Y(\u_ppwm/u_ex/_0303_ ),
    .A(net462),
    .B(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0863_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0291_ ),
    .A2(\u_ppwm/u_ex/_0293_ ),
    .Y(\u_ppwm/u_ex/_0304_ ),
    .B1(\u_ppwm/u_ex/_0292_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0864_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0303_ ),
    .A2(\u_ppwm/u_ex/_0304_ ),
    .Y(\u_ppwm/u_ex/_0305_ ),
    .B1(net358));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0865_  (.B1(\u_ppwm/u_ex/_0305_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0306_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0303_ ),
    .A2(\u_ppwm/u_ex/_0304_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0866_  (.A(net375),
    .B(net378),
    .C(\u_ppwm/u_ex/_0237_ ),
    .Y(\u_ppwm/u_ex/_0307_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0867_  (.A(\u_ppwm/u_ex/_0284_ ),
    .B(\u_ppwm/u_ex/_0307_ ),
    .Y(\u_ppwm/u_ex/_0308_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0868_  (.B1(\u_ppwm/u_ex/_0308_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0309_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0260_ ),
    .A2(\u_ppwm/u_ex/_0281_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0869_  (.A(\u_ppwm/pwm_value[7] ),
    .B(net385),
    .Y(\u_ppwm/u_ex/_0310_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0870_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0525_ ),
    .A2(net384),
    .Y(\u_ppwm/u_ex/_0311_ ),
    .B1(\u_ppwm/u_ex/_0310_ ));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0871_  (.A0(\u_ppwm/u_ex/_0286_ ),
    .A1(\u_ppwm/u_ex/_0311_ ),
    .S(net377),
    .X(\u_ppwm/u_ex/_0312_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0872_  (.Y(\u_ppwm/u_ex/_0313_ ),
    .B1(\u_ppwm/u_ex/_0312_ ),
    .B2(\u_ppwm/u_ex/_0240_ ),
    .A2(\u_ppwm/u_ex/_0256_ ),
    .A1(\u_ppwm/u_ex/_0233_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_ex/_0873_  (.A2(\u_ppwm/u_ex/_0313_ ),
    .A1(\u_ppwm/u_ex/_0309_ ),
    .B1(\u_ppwm/u_ex/_0232_ ),
    .X(\u_ppwm/u_ex/_0314_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0874_  (.Y(\u_ppwm/u_ex/_0315_ ),
    .B1(net365),
    .B2(\u_ppwm/global_counter[13] ),
    .A2(net367),
    .A1(\u_ppwm/global_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0875_  (.A(net360),
    .B(\u_ppwm/u_ex/_0315_ ),
    .Y(\u_ppwm/u_ex/_0316_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0876_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net450),
    .A2(\u_ppwm/u_ex/_0221_ ),
    .Y(\u_ppwm/u_ex/_0317_ ),
    .B1(\u_ppwm/u_ex/_0316_ ));
 sg13g2_nand4_1 \u_ppwm/u_ex/_0877_  (.B(\u_ppwm/u_ex/_0306_ ),
    .C(\u_ppwm/u_ex/_0314_ ),
    .A(\u_ppwm/u_ex/_0251_ ),
    .Y(\u_ppwm/u_ex/_0318_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0317_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0878_  (.B1(\u_ppwm/u_ex/_0318_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0319_ ),
    .VSS(VGND),
    .A1(net462),
    .A2(net354));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0879_  (.A(\u_ppwm/u_ex/_0032_ ),
    .B(\u_ppwm/u_ex/_0319_ ),
    .Y(\u_ppwm/u_ex/_0012_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0880_  (.Y(\u_ppwm/u_ex/_0320_ ),
    .A(net460),
    .B(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0881_  (.Y(\u_ppwm/u_ex/_0321_ ),
    .A(net460),
    .B(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0882_  (.A(\u_ppwm/u_ex/_0294_ ),
    .B(\u_ppwm/u_ex/_0303_ ),
    .Y(\u_ppwm/u_ex/_0322_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0883_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0029_ ),
    .A2(\u_ppwm/u_ex/_0030_ ),
    .Y(\u_ppwm/u_ex/_0323_ ),
    .B1(\u_ppwm/u_ex/_0035_ ));
 sg13g2_a21oi_2 \u_ppwm/u_ex/_0884_  (.VSS(VGND),
    .VDD(VPWR),
    .B1(\u_ppwm/u_ex/_0323_ ),
    .Y(\u_ppwm/u_ex/_0324_ ),
    .A2(\u_ppwm/u_ex/_0322_ ),
    .A1(\u_ppwm/u_ex/_0291_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0885_  (.B1(\u_ppwm/u_ex/_0224_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0325_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0321_ ),
    .A2(\u_ppwm/u_ex/_0324_ ));
 sg13g2_a21o_1 \u_ppwm/u_ex/_0886_  (.A2(\u_ppwm/u_ex/_0324_ ),
    .A1(\u_ppwm/u_ex/_0321_ ),
    .B1(\u_ppwm/u_ex/_0325_ ),
    .X(\u_ppwm/u_ex/_0326_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0887_  (.B1(\u_ppwm/u_ex/_0261_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0327_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0258_ ),
    .A2(\u_ppwm/u_ex/_0279_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0888_  (.Y(\u_ppwm/u_ex/_0328_ ),
    .B(net368),
    .A_N(\u_ppwm/u_ex/_0244_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0889_  (.B1(\u_ppwm/u_ex/_0328_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0329_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0239_ ),
    .A2(\u_ppwm/u_ex/_0281_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0890_  (.A(\u_ppwm/u_ex/_0327_ ),
    .B(\u_ppwm/u_ex/_0329_ ),
    .Y(\u_ppwm/u_ex/_0330_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0891_  (.A(net455),
    .B(net384),
    .Y(\u_ppwm/u_ex/_0331_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0892_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0524_ ),
    .A2(net384),
    .Y(\u_ppwm/u_ex/_0332_ ),
    .B1(\u_ppwm/u_ex/_0331_ ));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0893_  (.A0(\u_ppwm/u_ex/_0311_ ),
    .A1(\u_ppwm/u_ex/_0332_ ),
    .S(net377),
    .X(\u_ppwm/u_ex/_0333_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0894_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0241_ ),
    .C1(\u_ppwm/u_ex/_0330_ ),
    .B1(\u_ppwm/u_ex/_0333_ ),
    .A1(\u_ppwm/u_ex/_0234_ ),
    .Y(\u_ppwm/u_ex/_0334_ ),
    .A2(\u_ppwm/u_ex/_0288_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0895_  (.Y(\u_ppwm/u_ex/_0335_ ),
    .B1(net365),
    .B2(\u_ppwm/global_counter[14] ),
    .A2(net367),
    .A1(\u_ppwm/global_counter[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0896_  (.A(net359),
    .B(\u_ppwm/u_ex/_0335_ ),
    .Y(\u_ppwm/u_ex/_0336_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0897_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net449),
    .A2(\u_ppwm/u_ex/_0221_ ),
    .Y(\u_ppwm/u_ex/_0337_ ),
    .B1(\u_ppwm/u_ex/_0336_ ));
 sg13g2_nand4_1 \u_ppwm/u_ex/_0898_  (.B(\u_ppwm/u_ex/_0326_ ),
    .C(\u_ppwm/u_ex/_0334_ ),
    .A(net352),
    .Y(\u_ppwm/u_ex/_0338_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0337_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0899_  (.B1(net505),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0339_ ),
    .VSS(VGND),
    .A1(net460),
    .A2(net353));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0900_  (.A(\u_ppwm/u_ex/_0339_ ),
    .B_N(\u_ppwm/u_ex/_0338_ ),
    .Y(\u_ppwm/u_ex/_0013_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0901_  (.B1(\u_ppwm/u_ex/_0320_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0340_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0321_ ),
    .A2(\u_ppwm/u_ex/_0324_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0902_  (.B(net371),
    .A(net458),
    .X(\u_ppwm/u_ex/_0341_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0903_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0340_ ),
    .A2(\u_ppwm/u_ex/_0341_ ),
    .Y(\u_ppwm/u_ex/_0342_ ),
    .B1(net357));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0904_  (.B1(\u_ppwm/u_ex/_0342_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0343_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0340_ ),
    .A2(\u_ppwm/u_ex/_0341_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0905_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0236_ ),
    .A2(\u_ppwm/u_ex/_0278_ ),
    .Y(\u_ppwm/u_ex/_0344_ ),
    .B1(\u_ppwm/u_ex/_0262_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0906_  (.B1(\u_ppwm/u_ex/_0344_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0345_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0264_ ),
    .A2(\u_ppwm/u_ex/_0281_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0907_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net368),
    .A2(\u_ppwm/u_ex/_0243_ ),
    .Y(\u_ppwm/u_ex/_0346_ ),
    .B1(\u_ppwm/u_ex/_0345_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0908_  (.A(\u_ppwm/pwm_value[9] ),
    .B(net384),
    .Y(\u_ppwm/u_ex/_0347_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0909_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0523_ ),
    .A2(net384),
    .Y(\u_ppwm/u_ex/_0348_ ),
    .B1(\u_ppwm/u_ex/_0347_ ));
 sg13g2_mux2_1 \u_ppwm/u_ex/_0910_  (.A0(\u_ppwm/u_ex/_0332_ ),
    .A1(\u_ppwm/u_ex/_0348_ ),
    .S(net377),
    .X(\u_ppwm/u_ex/_0349_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0911_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0241_ ),
    .C1(\u_ppwm/u_ex/_0346_ ),
    .B1(\u_ppwm/u_ex/_0349_ ),
    .A1(\u_ppwm/u_ex/_0234_ ),
    .Y(\u_ppwm/u_ex/_0350_ ),
    .A2(\u_ppwm/u_ex/_0312_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0912_  (.Y(\u_ppwm/u_ex/_0351_ ),
    .B1(net365),
    .B2(\u_ppwm/global_counter[15] ),
    .A2(net367),
    .A1(\u_ppwm/global_counter[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0913_  (.A(net359),
    .B(\u_ppwm/u_ex/_0351_ ),
    .Y(\u_ppwm/u_ex/_0352_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0914_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/reg_value_q[5] ),
    .A2(\u_ppwm/u_ex/_0221_ ),
    .Y(\u_ppwm/u_ex/_0353_ ),
    .B1(\u_ppwm/u_ex/_0352_ ));
 sg13g2_nand4_1 \u_ppwm/u_ex/_0915_  (.B(\u_ppwm/u_ex/_0343_ ),
    .C(\u_ppwm/u_ex/_0350_ ),
    .A(net353),
    .Y(\u_ppwm/u_ex/_0354_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0353_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0916_  (.B1(net491),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0355_ ),
    .VSS(VGND),
    .A1(net458),
    .A2(net352));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0917_  (.A(\u_ppwm/u_ex/_0355_ ),
    .B_N(\u_ppwm/u_ex/_0354_ ),
    .Y(\u_ppwm/u_ex/_0014_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0918_  (.A(net456),
    .B(net371),
    .Y(\u_ppwm/u_ex/_0356_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_ex/_0919_  (.A(net456),
    .B(net371),
    .X(\u_ppwm/u_ex/_0357_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0920_  (.A(\u_ppwm/u_ex/_0356_ ),
    .B(\u_ppwm/u_ex/_0357_ ),
    .Y(\u_ppwm/u_ex/_0358_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0921_  (.B1(net371),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0359_ ),
    .VSS(VGND),
    .A1(net458),
    .A2(net460));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_0922_  (.Y(\u_ppwm/u_ex/_0360_ ),
    .B(\u_ppwm/u_ex/_0341_ ),
    .A_N(\u_ppwm/u_ex/_0321_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0923_  (.B1(\u_ppwm/u_ex/_0359_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0361_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0324_ ),
    .A2(\u_ppwm/u_ex/_0360_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0924_  (.B(\u_ppwm/u_ex/_0361_ ),
    .A(\u_ppwm/u_ex/_0358_ ),
    .X(\u_ppwm/u_ex/_0362_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0925_  (.Y(\u_ppwm/u_ex/_0363_ ),
    .A(net368),
    .B(\u_ppwm/u_ex/_0254_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0926_  (.Y(\u_ppwm/u_ex/_0364_ ),
    .B1(\u_ppwm/u_ex/_0280_ ),
    .B2(\u_ppwm/u_ex/_0245_ ),
    .A2(\u_ppwm/u_ex/_0278_ ),
    .A1(\u_ppwm/u_ex/_0237_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0927_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0363_ ),
    .A2(\u_ppwm/u_ex/_0364_ ),
    .Y(\u_ppwm/u_ex/_0365_ ),
    .B1(\u_ppwm/u_ex/_0262_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_0928_  (.A(net370),
    .B(\u_ppwm/u_ex/_0348_ ),
    .X(\u_ppwm/u_ex/_0366_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0929_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_ex/_0241_ ),
    .C1(\u_ppwm/u_ex/_0365_ ),
    .B1(\u_ppwm/u_ex/_0366_ ),
    .A1(\u_ppwm/u_ex/_0234_ ),
    .Y(\u_ppwm/u_ex/_0367_ ),
    .A2(\u_ppwm/u_ex/_0333_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0930_  (.Y(\u_ppwm/u_ex/_0368_ ),
    .B1(net365),
    .B2(net439),
    .A2(net367),
    .A1(\u_ppwm/global_counter[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0931_  (.A(net361),
    .B(\u_ppwm/u_ex/_0368_ ),
    .Y(\u_ppwm/u_ex/_0369_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0932_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net448),
    .A2(\u_ppwm/u_ex/_0221_ ),
    .Y(\u_ppwm/u_ex/_0370_ ),
    .B1(\u_ppwm/u_ex/_0369_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_0933_  (.B(\u_ppwm/u_ex/_0367_ ),
    .C(\u_ppwm/u_ex/_0370_ ),
    .A(net352),
    .Y(\u_ppwm/u_ex/_0371_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0934_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0224_ ),
    .A2(\u_ppwm/u_ex/_0362_ ),
    .Y(\u_ppwm/u_ex/_0372_ ),
    .B1(\u_ppwm/u_ex/_0371_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0935_  (.B1(net491),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0373_ ),
    .VSS(VGND),
    .A1(net456),
    .A2(net352));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0936_  (.A(\u_ppwm/u_ex/_0372_ ),
    .B(\u_ppwm/u_ex/_0373_ ),
    .Y(\u_ppwm/u_ex/_0015_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0937_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0358_ ),
    .A2(\u_ppwm/u_ex/_0361_ ),
    .Y(\u_ppwm/u_ex/_0374_ ),
    .B1(\u_ppwm/u_ex/_0357_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0938_  (.Y(\u_ppwm/u_ex/_0375_ ),
    .A(net664),
    .B(net371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0939_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0374_ ),
    .A2(\u_ppwm/u_ex/_0375_ ),
    .Y(\u_ppwm/u_ex/_0376_ ),
    .B1(net357));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0940_  (.B1(\u_ppwm/u_ex/_0376_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0377_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0374_ ),
    .A2(\u_ppwm/u_ex/_0375_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0941_  (.Y(\u_ppwm/u_ex/_0378_ ),
    .B1(\u_ppwm/u_ex/_0286_ ),
    .B2(net368),
    .A2(\u_ppwm/u_ex/_0278_ ),
    .A1(\u_ppwm/u_ex/_0244_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0942_  (.B1(\u_ppwm/u_ex/_0378_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0379_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0257_ ),
    .A2(\u_ppwm/u_ex/_0281_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0943_  (.Y(\u_ppwm/u_ex/_0380_ ),
    .B1(\u_ppwm/u_ex/_0379_ ),
    .B2(\u_ppwm/u_ex/_0261_ ),
    .A2(\u_ppwm/u_ex/_0349_ ),
    .A1(\u_ppwm/u_ex/_0234_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0944_  (.B1(\u_ppwm/u_ex/reg_value_q[7] ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0381_ ),
    .VSS(VGND),
    .A1(net381),
    .A2(net370));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0945_  (.Y(\u_ppwm/u_ex/_0382_ ),
    .B1(net364),
    .B2(\u_ppwm/global_counter[17] ),
    .A2(net366),
    .A1(\u_ppwm/global_counter[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_ex/_0946_  (.A2(\u_ppwm/u_ex/_0382_ ),
    .A1(\u_ppwm/u_ex/_0381_ ),
    .B1(net361),
    .X(\u_ppwm/u_ex/_0383_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 \u_ppwm/u_ex/_0947_  (.X(\u_ppwm/u_ex/_0384_ ),
    .A(net352),
    .B(\u_ppwm/u_ex/_0380_ ),
    .C(\u_ppwm/u_ex/_0383_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0948_  (.B1(net491),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0385_ ),
    .VSS(VGND),
    .A1(net664),
    .A2(net352));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0949_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0377_ ),
    .A2(\u_ppwm/u_ex/_0384_ ),
    .Y(\u_ppwm/u_ex/_0016_ ),
    .B1(\u_ppwm/u_ex/_0385_ ));
 sg13g2_or4_1 \u_ppwm/u_ex/_0950_  (.A(\u_ppwm/u_ex/_0356_ ),
    .B(\u_ppwm/u_ex/_0357_ ),
    .C(\u_ppwm/u_ex/_0360_ ),
    .D(\u_ppwm/u_ex/_0375_ ),
    .X(\u_ppwm/u_ex/_0386_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0951_  (.B1(net371),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0387_ ),
    .VSS(VGND),
    .A1(\u_ppwm/pwm_value[7] ),
    .A2(net456));
 sg13g2_and2_1 \u_ppwm/u_ex/_0952_  (.A(\u_ppwm/u_ex/_0359_ ),
    .B(\u_ppwm/u_ex/_0387_ ),
    .X(\u_ppwm/u_ex/_0388_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0953_  (.B1(\u_ppwm/u_ex/_0388_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0389_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0324_ ),
    .A2(\u_ppwm/u_ex/_0386_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0954_  (.A(\u_ppwm/u_ex/_0531_ ),
    .B(\u_ppwm/u_ex/_0035_ ),
    .Y(\u_ppwm/u_ex/_0390_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0955_  (.B(net372),
    .A(net455),
    .X(\u_ppwm/u_ex/_0391_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0956_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0389_ ),
    .A2(\u_ppwm/u_ex/_0391_ ),
    .Y(\u_ppwm/u_ex/_0392_ ),
    .B1(net357));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0957_  (.B1(\u_ppwm/u_ex/_0392_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0393_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0389_ ),
    .A2(\u_ppwm/u_ex/_0391_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0958_  (.Y(\u_ppwm/u_ex/_0394_ ),
    .B1(\u_ppwm/u_ex/_0311_ ),
    .B2(net368),
    .A2(\u_ppwm/u_ex/_0278_ ),
    .A1(\u_ppwm/u_ex/_0242_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0959_  (.B1(\u_ppwm/u_ex/_0394_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0395_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0281_ ),
    .A2(\u_ppwm/u_ex/_0289_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0960_  (.Y(\u_ppwm/u_ex/_0396_ ),
    .B1(\u_ppwm/u_ex/_0395_ ),
    .B2(\u_ppwm/u_ex/_0261_ ),
    .A2(\u_ppwm/u_ex/_0366_ ),
    .A1(\u_ppwm/u_ex/_0234_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0961_  (.Y(\u_ppwm/u_ex/_0397_ ),
    .B1(net364),
    .B2(\u_ppwm/global_counter[18] ),
    .A2(net366),
    .A1(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0962_  (.A(net361),
    .B(\u_ppwm/u_ex/_0397_ ),
    .Y(\u_ppwm/u_ex/_0398_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0963_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net663),
    .A2(\u_ppwm/u_ex/_0221_ ),
    .Y(\u_ppwm/u_ex/_0399_ ),
    .B1(\u_ppwm/u_ex/_0398_ ));
 sg13g2_nand4_1 \u_ppwm/u_ex/_0964_  (.B(\u_ppwm/u_ex/_0393_ ),
    .C(\u_ppwm/u_ex/_0396_ ),
    .A(net352),
    .Y(\u_ppwm/u_ex/_0400_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0399_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0965_  (.B1(net490),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0401_ ),
    .VSS(VGND),
    .A1(net455),
    .A2(net352));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0966_  (.A(\u_ppwm/u_ex/_0401_ ),
    .B_N(\u_ppwm/u_ex/_0400_ ),
    .Y(\u_ppwm/u_ex/_0017_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0967_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0389_ ),
    .A2(\u_ppwm/u_ex/_0391_ ),
    .Y(\u_ppwm/u_ex/_0402_ ),
    .B1(\u_ppwm/u_ex/_0390_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0968_  (.Y(\u_ppwm/u_ex/_0403_ ),
    .A(net454),
    .B(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0969_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0402_ ),
    .A2(\u_ppwm/u_ex/_0403_ ),
    .Y(\u_ppwm/u_ex/_0404_ ),
    .B1(net357));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0970_  (.B1(\u_ppwm/u_ex/_0404_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0405_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0402_ ),
    .A2(\u_ppwm/u_ex/_0403_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0971_  (.Y(\u_ppwm/u_ex/_0406_ ),
    .B1(\u_ppwm/u_ex/_0332_ ),
    .B2(net368),
    .A2(\u_ppwm/u_ex/_0312_ ),
    .A1(\u_ppwm/u_ex/_0280_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0972_  (.B1(\u_ppwm/u_ex/_0406_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0407_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0255_ ),
    .A2(\u_ppwm/u_ex/_0279_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_0973_  (.A(\u_ppwm/u_ex/_0523_ ),
    .B(net366),
    .C(net364),
    .Y(\u_ppwm/u_ex/_0408_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_0974_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/global_counter[19] ),
    .C1(\u_ppwm/u_ex/_0408_ ),
    .B1(net364),
    .A1(net441),
    .Y(\u_ppwm/u_ex/_0409_ ),
    .A2(net366));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0975_  (.B1(net353),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0410_ ),
    .VSS(VGND),
    .A1(net361),
    .A2(\u_ppwm/u_ex/_0409_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0976_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0261_ ),
    .A2(\u_ppwm/u_ex/_0407_ ),
    .Y(\u_ppwm/u_ex/_0411_ ),
    .B1(\u_ppwm/u_ex/_0410_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0977_  (.B1(net492),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0412_ ),
    .VSS(VGND),
    .A1(net454),
    .A2(net353));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0978_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0405_ ),
    .A2(\u_ppwm/u_ex/_0411_ ),
    .Y(\u_ppwm/u_ex/_0018_ ),
    .B1(\u_ppwm/u_ex/_0412_ ));
 sg13g2_nor2_2 \u_ppwm/u_ex/_0979_  (.A(\u_ppwm/u_ex/_0034_ ),
    .B(net363),
    .Y(\u_ppwm/u_ex/_0413_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0980_  (.Y(\u_ppwm/u_ex/_0414_ ),
    .A(\u_ppwm/global_counter[10] ),
    .B(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0981_  (.Y(\u_ppwm/u_ex/_0415_ ),
    .B1(net356),
    .B2(net445),
    .A2(net362),
    .A1(\u_ppwm/pwm_value[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_ex/_0982_  (.A2(\u_ppwm/u_ex/_0415_ ),
    .A1(\u_ppwm/u_ex/_0414_ ),
    .B1(net360),
    .X(\u_ppwm/u_ex/_0416_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0983_  (.A(net379),
    .B(\u_ppwm/u_ex/_0135_ ),
    .Y(\u_ppwm/u_ex/_0417_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0984_  (.Y(\u_ppwm/u_ex/_0418_ ),
    .B1(\u_ppwm/u_ex/_0417_ ),
    .B2(\u_ppwm/u_ex/_0219_ ),
    .A2(\u_ppwm/u_ex/_0248_ ),
    .A1(net385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_0985_  (.A(\u_ppwm/u_ex/_0418_ ),
    .B_N(net446),
    .Y(\u_ppwm/u_ex/_0419_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_ex/_0986_  (.A(\u_ppwm/u_ex/reg_value_q[0] ),
    .B(net383),
    .X(\u_ppwm/u_ex/_0420_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0987_  (.B(\u_ppwm/instr[4] ),
    .A(\u_ppwm/u_ex/reg_value_q[0] ),
    .X(\u_ppwm/u_ex/_0421_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0988_  (.Y(\u_ppwm/u_ex/_0422_ ),
    .B1(\u_ppwm/u_ex/_0421_ ),
    .B2(\u_ppwm/u_ex/_0224_ ),
    .A2(\u_ppwm/u_ex/_0228_ ),
    .A1(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_ex/_0989_  (.B(\u_ppwm/u_ex/_0416_ ),
    .C(net350),
    .A(\u_ppwm/u_ex/_0246_ ),
    .Y(\u_ppwm/u_ex/_0423_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0422_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_0990_  (.B1(\u_ppwm/u_ex/_0423_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0424_ ),
    .VSS(VGND),
    .A1(net660),
    .A2(net350));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0991_  (.A(\u_ppwm/u_ex/_0032_ ),
    .B(\u_ppwm/u_ex/_0424_ ),
    .Y(\u_ppwm/u_ex/_0019_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_ex/_0992_  (.A(net453),
    .B(net380),
    .X(\u_ppwm/u_ex/_0425_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_0993_  (.B(net380),
    .A(net453),
    .X(\u_ppwm/u_ex/_0426_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_0994_  (.Y(\u_ppwm/u_ex/_0427_ ),
    .A(\u_ppwm/u_ex/_0420_ ),
    .B(\u_ppwm/u_ex/_0426_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_0995_  (.A(net358),
    .B(\u_ppwm/u_ex/_0427_ ),
    .Y(\u_ppwm/u_ex/_0428_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0996_  (.Y(\u_ppwm/u_ex/_0429_ ),
    .A(\u_ppwm/u_ex/_0267_ ),
    .B(net350),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_0997_  (.Y(\u_ppwm/u_ex/_0430_ ),
    .A(net444),
    .B(net356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_0998_  (.Y(\u_ppwm/u_ex/_0431_ ),
    .B1(net355),
    .B2(\u_ppwm/global_counter[11] ),
    .A2(net362),
    .A1(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_0999_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0430_ ),
    .A2(\u_ppwm/u_ex/_0431_ ),
    .Y(\u_ppwm/u_ex/_0432_ ),
    .B1(net360));
 sg13g2_nor4_1 \u_ppwm/u_ex/_1000_  (.A(\u_ppwm/u_ex/_0266_ ),
    .B(\u_ppwm/u_ex/_0428_ ),
    .C(\u_ppwm/u_ex/_0429_ ),
    .D(\u_ppwm/u_ex/_0432_ ),
    .Y(\u_ppwm/u_ex/_0433_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1001_  (.B1(net506),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0434_ ),
    .VSS(VGND),
    .A1(net453),
    .A2(net350));
 sg13g2_nor2_1 \u_ppwm/u_ex/_1002_  (.A(\u_ppwm/u_ex/_0433_ ),
    .B(\u_ppwm/u_ex/_0434_ ),
    .Y(\u_ppwm/u_ex/_0020_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1003_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0420_ ),
    .A2(\u_ppwm/u_ex/_0426_ ),
    .Y(\u_ppwm/u_ex/_0435_ ),
    .B1(\u_ppwm/u_ex/_0425_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1004_  (.Y(\u_ppwm/u_ex/_0436_ ),
    .A(net451),
    .B(net376),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_1005_  (.Y(\u_ppwm/u_ex/_0437_ ),
    .A(net451),
    .B(net376),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 \u_ppwm/u_ex/_1006_  (.VSS(VGND),
    .VDD(VPWR),
    .X(\u_ppwm/u_ex/_0438_ ),
    .B(\u_ppwm/u_ex/_0437_ ),
    .A(\u_ppwm/u_ex/_0435_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1007_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0435_ ),
    .A2(\u_ppwm/u_ex/_0437_ ),
    .Y(\u_ppwm/u_ex/_0439_ ),
    .B1(net358));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1008_  (.Y(\u_ppwm/u_ex/_0440_ ),
    .A(net443),
    .B(\u_ppwm/u_ex/_0188_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_1009_  (.Y(\u_ppwm/u_ex/_0441_ ),
    .B1(net355),
    .B2(net440),
    .A2(net362),
    .A1(\u_ppwm/pwm_value[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1010_  (.Y(\u_ppwm/u_ex/_0442_ ),
    .A(\u_ppwm/u_ex/_0440_ ),
    .B(\u_ppwm/u_ex/_0441_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_1011_  (.Y(\u_ppwm/u_ex/_0443_ ),
    .B1(\u_ppwm/u_ex/_0442_ ),
    .B2(\u_ppwm/u_ex/_0219_ ),
    .A2(\u_ppwm/u_ex/_0439_ ),
    .A1(\u_ppwm/u_ex/_0438_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_ex/_1012_  (.B(\u_ppwm/u_ex/_0298_ ),
    .C(net350),
    .A(\u_ppwm/u_ex/_0290_ ),
    .Y(\u_ppwm/u_ex/_0444_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0443_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1013_  (.B1(net508),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0445_ ),
    .VSS(VGND),
    .A1(net451),
    .A2(net350));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_1014_  (.A(\u_ppwm/u_ex/_0445_ ),
    .B_N(\u_ppwm/u_ex/_0444_ ),
    .Y(\u_ppwm/u_ex/_0021_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_1015_  (.Y(\u_ppwm/u_ex/_0446_ ),
    .A(net450),
    .B(net376),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1016_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0436_ ),
    .A2(\u_ppwm/u_ex/_0438_ ),
    .Y(\u_ppwm/u_ex/_0447_ ),
    .B1(\u_ppwm/u_ex/_0446_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_1017_  (.B(\u_ppwm/u_ex/_0438_ ),
    .C(\u_ppwm/u_ex/_0446_ ),
    .A(\u_ppwm/u_ex/_0436_ ),
    .Y(\u_ppwm/u_ex/_0448_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_1018_  (.A(net358),
    .B(\u_ppwm/u_ex/_0447_ ),
    .Y(\u_ppwm/u_ex/_0449_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_ex/_1019_  (.A(net387),
    .B(\u_ppwm/u_ex/_0043_ ),
    .C(net362),
    .Y(\u_ppwm/u_ex/_0450_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_1020_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/global_counter[13] ),
    .C1(\u_ppwm/u_ex/_0450_ ),
    .B1(net355),
    .A1(net692),
    .Y(\u_ppwm/u_ex/_0451_ ),
    .A2(net362));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1021_  (.B1(net351),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0452_ ),
    .VSS(VGND),
    .A1(net360),
    .A2(\u_ppwm/u_ex/_0451_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1022_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0448_ ),
    .A2(\u_ppwm/u_ex/_0449_ ),
    .Y(\u_ppwm/u_ex/_0453_ ),
    .B1(\u_ppwm/u_ex/_0452_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1023_  (.B1(net506),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0454_ ),
    .VSS(VGND),
    .A1(net450),
    .A2(net350));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1024_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0314_ ),
    .A2(\u_ppwm/u_ex/_0453_ ),
    .Y(\u_ppwm/u_ex/_0022_ ),
    .B1(\u_ppwm/u_ex/_0454_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_1025_  (.A(\u_ppwm/u_ex/_0528_ ),
    .B(\u_ppwm/u_ex/_0035_ ),
    .Y(\u_ppwm/u_ex/_0455_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_1026_  (.B(net373),
    .A(net449),
    .X(\u_ppwm/u_ex/_0456_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 \u_ppwm/u_ex/_1027_  (.VSS(VGND),
    .VDD(VPWR),
    .X(\u_ppwm/u_ex/_0457_ ),
    .B(\u_ppwm/u_ex/_0446_ ),
    .A(\u_ppwm/u_ex/_0437_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1028_  (.B1(net376),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0458_ ),
    .VSS(VGND),
    .A1(net450),
    .A2(net451));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1029_  (.B1(\u_ppwm/u_ex/_0458_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0459_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0435_ ),
    .A2(\u_ppwm/u_ex/_0457_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1030_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0456_ ),
    .A2(\u_ppwm/u_ex/_0459_ ),
    .Y(\u_ppwm/u_ex/_0460_ ),
    .B1(net357));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1031_  (.B1(\u_ppwm/u_ex/_0460_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0461_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0456_ ),
    .A2(\u_ppwm/u_ex/_0459_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1032_  (.Y(\u_ppwm/u_ex/_0462_ ),
    .A(\u_ppwm/global_counter[4] ),
    .B(net356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_1033_  (.Y(\u_ppwm/u_ex/_0463_ ),
    .B1(net355),
    .B2(\u_ppwm/global_counter[14] ),
    .A2(net362),
    .A1(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_ex/_1034_  (.A2(\u_ppwm/u_ex/_0463_ ),
    .A1(\u_ppwm/u_ex/_0462_ ),
    .B1(net359),
    .X(\u_ppwm/u_ex/_0464_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_ex/_1035_  (.B(net351),
    .C(\u_ppwm/u_ex/_0461_ ),
    .A(\u_ppwm/u_ex/_0334_ ),
    .Y(\u_ppwm/u_ex/_0465_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0464_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1036_  (.B1(net505),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0466_ ),
    .VSS(VGND),
    .A1(net449),
    .A2(net349));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_1037_  (.A(\u_ppwm/u_ex/_0466_ ),
    .B_N(\u_ppwm/u_ex/_0465_ ),
    .Y(\u_ppwm/u_ex/_0023_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1038_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0456_ ),
    .A2(\u_ppwm/u_ex/_0459_ ),
    .Y(\u_ppwm/u_ex/_0467_ ),
    .B1(\u_ppwm/u_ex/_0455_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_1039_  (.B(net373),
    .A(\u_ppwm/u_ex/reg_value_q[5] ),
    .X(\u_ppwm/u_ex/_0468_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_1040_  (.Y(\u_ppwm/u_ex/_0469_ ),
    .A(\u_ppwm/u_ex/reg_value_q[5] ),
    .B(net373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1041_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0467_ ),
    .A2(\u_ppwm/u_ex/_0469_ ),
    .Y(\u_ppwm/u_ex/_0470_ ),
    .B1(net358));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1042_  (.B1(\u_ppwm/u_ex/_0470_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0471_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0467_ ),
    .A2(\u_ppwm/u_ex/_0469_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1043_  (.Y(\u_ppwm/u_ex/_0472_ ),
    .A(\u_ppwm/global_counter[15] ),
    .B(\u_ppwm/u_ex/_0413_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_1044_  (.Y(\u_ppwm/u_ex/_0473_ ),
    .B1(\u_ppwm/u_ex/_0188_ ),
    .B2(\u_ppwm/global_counter[5] ),
    .A2(net362),
    .A1(net459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_ex/_1045_  (.A2(\u_ppwm/u_ex/_0473_ ),
    .A1(\u_ppwm/u_ex/_0472_ ),
    .B1(net359),
    .X(\u_ppwm/u_ex/_0474_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_ex/_1046_  (.B(net351),
    .C(\u_ppwm/u_ex/_0471_ ),
    .A(\u_ppwm/u_ex/_0350_ ),
    .Y(\u_ppwm/u_ex/_0475_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0474_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1047_  (.B1(net506),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0476_ ),
    .VSS(VGND),
    .A1(net667),
    .A2(net351));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_1048_  (.A(\u_ppwm/u_ex/_0476_ ),
    .B_N(\u_ppwm/u_ex/_0475_ ),
    .Y(\u_ppwm/u_ex/_0024_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_1049_  (.A(\u_ppwm/u_ex/_0526_ ),
    .B(\u_ppwm/u_ex/_0035_ ),
    .Y(\u_ppwm/u_ex/_0477_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_ex/_1050_  (.B(net373),
    .A(net448),
    .X(\u_ppwm/u_ex/_0478_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_ex/_1051_  (.VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0479_ ),
    .A(\u_ppwm/u_ex/_0478_ ),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1052_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0527_ ),
    .A2(\u_ppwm/u_ex/_0528_ ),
    .Y(\u_ppwm/u_ex/_0480_ ),
    .B1(\u_ppwm/u_ex/_0035_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_1053_  (.A(\u_ppwm/u_ex/_0456_ ),
    .B(\u_ppwm/u_ex/_0468_ ),
    .X(\u_ppwm/u_ex/_0481_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1054_  (.Y(\u_ppwm/u_ex/_0482_ ),
    .A(\u_ppwm/u_ex/_0456_ ),
    .B(\u_ppwm/u_ex/_0468_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_ex/_1055_  (.A2(\u_ppwm/u_ex/_0481_ ),
    .A1(\u_ppwm/u_ex/_0459_ ),
    .B1(\u_ppwm/u_ex/_0480_ ),
    .X(\u_ppwm/u_ex/_0483_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1056_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0478_ ),
    .A2(\u_ppwm/u_ex/_0483_ ),
    .Y(\u_ppwm/u_ex/_0484_ ),
    .B1(net357));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1057_  (.B1(\u_ppwm/u_ex/_0484_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0485_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0478_ ),
    .A2(\u_ppwm/u_ex/_0483_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1058_  (.Y(\u_ppwm/u_ex/_0486_ ),
    .A(\u_ppwm/global_counter[6] ),
    .B(net356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_1059_  (.Y(\u_ppwm/u_ex/_0487_ ),
    .B1(\u_ppwm/u_ex/_0413_ ),
    .B2(\u_ppwm/global_counter[16] ),
    .A2(net362),
    .A1(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_ex/_1060_  (.A2(\u_ppwm/u_ex/_0487_ ),
    .A1(\u_ppwm/u_ex/_0486_ ),
    .B1(net359),
    .X(\u_ppwm/u_ex/_0488_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_ex/_1061_  (.B(net349),
    .C(\u_ppwm/u_ex/_0485_ ),
    .A(\u_ppwm/u_ex/_0367_ ),
    .Y(\u_ppwm/u_ex/_0489_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0488_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1062_  (.B1(net505),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0490_ ),
    .VSS(VGND),
    .A1(net448),
    .A2(net349));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_1063_  (.A(\u_ppwm/u_ex/_0490_ ),
    .B_N(\u_ppwm/u_ex/_0489_ ),
    .Y(\u_ppwm/u_ex/_0025_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1064_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0478_ ),
    .A2(\u_ppwm/u_ex/_0483_ ),
    .Y(\u_ppwm/u_ex/_0491_ ),
    .B1(\u_ppwm/u_ex/_0477_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_1065_  (.Y(\u_ppwm/u_ex/_0492_ ),
    .A(net662),
    .B(net373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1066_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0491_ ),
    .A2(\u_ppwm/u_ex/_0492_ ),
    .Y(\u_ppwm/u_ex/_0493_ ),
    .B1(net358));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1067_  (.B1(\u_ppwm/u_ex/_0493_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0494_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0491_ ),
    .A2(\u_ppwm/u_ex/_0492_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1068_  (.Y(\u_ppwm/u_ex/_0495_ ),
    .A(net645),
    .B(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_1069_  (.Y(\u_ppwm/u_ex/_0496_ ),
    .B1(net356),
    .B2(net630),
    .A2(net363),
    .A1(\u_ppwm/pwm_value[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1070_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0495_ ),
    .A2(\u_ppwm/u_ex/_0496_ ),
    .Y(\u_ppwm/u_ex/_0497_ ),
    .B1(net361));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1071_  (.Y(\u_ppwm/u_ex/_0498_ ),
    .A(\u_ppwm/u_ex/_0380_ ),
    .B(net349),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_ex/_1072_  (.A(\u_ppwm/u_ex/_0497_ ),
    .B(\u_ppwm/u_ex/_0498_ ),
    .Y(\u_ppwm/u_ex/_0499_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1073_  (.B1(net505),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0500_ ),
    .VSS(VGND),
    .A1(net662),
    .A2(net349));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1074_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0494_ ),
    .A2(\u_ppwm/u_ex/_0499_ ),
    .Y(\u_ppwm/u_ex/_0026_ ),
    .B1(\u_ppwm/u_ex/_0500_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_1075_  (.A(\u_ppwm/u_ex/_0479_ ),
    .B(\u_ppwm/u_ex/_0482_ ),
    .C(\u_ppwm/u_ex/_0492_ ),
    .Y(\u_ppwm/u_ex/_0501_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1076_  (.B1(net373),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0502_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/reg_value_q[7] ),
    .A2(net448));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_1077_  (.Y(\u_ppwm/u_ex/_0503_ ),
    .B(\u_ppwm/u_ex/_0502_ ),
    .A_N(\u_ppwm/u_ex/_0480_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 \u_ppwm/u_ex/_1078_  (.VSS(VGND),
    .VDD(VPWR),
    .B1(\u_ppwm/u_ex/_0503_ ),
    .Y(\u_ppwm/u_ex/_0504_ ),
    .A2(\u_ppwm/u_ex/_0501_ ),
    .A1(\u_ppwm/u_ex/_0459_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1079_  (.Y(\u_ppwm/u_ex/_0505_ ),
    .A(\u_ppwm/u_ex/reg_value_q[8] ),
    .B(net371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_1080_  (.Y(\u_ppwm/u_ex/_0506_ ),
    .A(\u_ppwm/u_ex/reg_value_q[8] ),
    .B(net371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1081_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0504_ ),
    .A2(\u_ppwm/u_ex/_0506_ ),
    .Y(\u_ppwm/u_ex/_0507_ ),
    .B1(net357));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1082_  (.B1(\u_ppwm/u_ex/_0507_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0508_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0504_ ),
    .A2(\u_ppwm/u_ex/_0506_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_1083_  (.Y(\u_ppwm/u_ex/_0509_ ),
    .A(\u_ppwm/global_counter[18] ),
    .B(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_1084_  (.Y(\u_ppwm/u_ex/_0510_ ),
    .B1(net356),
    .B2(net442),
    .A2(net363),
    .A1(\u_ppwm/pwm_value[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_ex/_1085_  (.A2(\u_ppwm/u_ex/_0510_ ),
    .A1(\u_ppwm/u_ex/_0509_ ),
    .B1(net361),
    .X(\u_ppwm/u_ex/_0511_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_ex/_1086_  (.B(net349),
    .C(\u_ppwm/u_ex/_0508_ ),
    .A(\u_ppwm/u_ex/_0396_ ),
    .Y(\u_ppwm/u_ex/_0512_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_ex/_0511_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1087_  (.B1(net491),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0513_ ),
    .VSS(VGND),
    .A1(net663),
    .A2(net349));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_1088_  (.A(\u_ppwm/u_ex/_0513_ ),
    .B_N(\u_ppwm/u_ex/_0512_ ),
    .Y(\u_ppwm/u_ex/_0027_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1089_  (.B1(\u_ppwm/u_ex/_0505_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0514_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0504_ ),
    .A2(\u_ppwm/u_ex/_0506_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_1090_  (.B(net374),
    .A(net657),
    .X(\u_ppwm/u_ex/_0515_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1091_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0514_ ),
    .A2(\u_ppwm/u_ex/_0515_ ),
    .Y(\u_ppwm/u_ex/_0516_ ),
    .B1(net357));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1092_  (.B1(\u_ppwm/u_ex/_0516_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0517_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_ex/_0514_ ),
    .A2(\u_ppwm/u_ex/_0515_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1093_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net381),
    .A2(net370),
    .Y(\u_ppwm/u_ex/_0518_ ),
    .B1(\u_ppwm/u_ex/_0530_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_1094_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/global_counter[19] ),
    .C1(\u_ppwm/u_ex/_0518_ ),
    .B1(net355),
    .A1(net441),
    .Y(\u_ppwm/u_ex/_0519_ ),
    .A2(net356));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1095_  (.B1(net350),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0520_ ),
    .VSS(VGND),
    .A1(net361),
    .A2(\u_ppwm/u_ex/_0519_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1096_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0261_ ),
    .A2(\u_ppwm/u_ex/_0407_ ),
    .Y(\u_ppwm/u_ex/_0521_ ),
    .B1(\u_ppwm/u_ex/_0520_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_1097_  (.B1(net491),
    .VDD(VPWR),
    .Y(\u_ppwm/u_ex/_0522_ ),
    .VSS(VGND),
    .A1(net657),
    .A2(net349));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_1098_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_ex/_0517_ ),
    .A2(\u_ppwm/u_ex/_0521_ ),
    .Y(\u_ppwm/u_ex/_0028_ ),
    .B1(\u_ppwm/u_ex/_0522_ ));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1099_  (.RESET_B(net52),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0003_ ),
    .Q(\u_ppwm/pc[0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1100_  (.RESET_B(net51),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0004_ ),
    .Q(\u_ppwm/pc[1] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1101_  (.RESET_B(net49),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0005_ ),
    .Q(\u_ppwm/pc[2] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1102_  (.RESET_B(net47),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net685),
    .Q(\u_ppwm/pc[3] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1103_  (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net650),
    .Q(\u_ppwm/u_ex/cmp_flag_q ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1104_  (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net248),
    .Q(\u_ppwm/polarity ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1105_  (.RESET_B(net41),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net661),
    .Q(\u_ppwm/pwm_value[0] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1106_  (.RESET_B(net39),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net688),
    .Q(\u_ppwm/pwm_value[1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1107_  (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0011_ ),
    .Q(\u_ppwm/pwm_value[2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1108_  (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0012_ ),
    .Q(\u_ppwm/pwm_value[3] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1109_  (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0013_ ),
    .Q(\u_ppwm/pwm_value[4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1110_  (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net670),
    .Q(\u_ppwm/pwm_value[5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1111_  (.RESET_B(net29),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0015_ ),
    .Q(\u_ppwm/pwm_value[6] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1112_  (.RESET_B(net27),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0016_ ),
    .Q(\u_ppwm/pwm_value[7] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1113_  (.RESET_B(net50),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0017_ ),
    .Q(\u_ppwm/pwm_value[8] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1114_  (.RESET_B(net46),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0018_ ),
    .Q(\u_ppwm/pwm_value[9] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1115_  (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0019_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1116_  (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net679),
    .Q(\u_ppwm/u_ex/reg_value_q[1] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1117_  (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0021_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1118_  (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0022_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[3] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1119_  (.RESET_B(net26),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0023_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1120_  (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0024_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[5] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1121_  (.RESET_B(net36),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0025_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[6] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1122_  (.RESET_B(net28),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0026_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1123_  (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_ex/_0027_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[8] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_1124_  (.RESET_B(net53),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net658),
    .Q(\u_ppwm/u_ex/reg_value_q[9] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1125_  (.RESET_B(net54),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net616),
    .Q(\u_ppwm/u_ex/state_q[0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1126_  (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net219),
    .Q(\u_ppwm/u_ex/state_q[1] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_1127_  (.RESET_B(net48),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net643),
    .Q(\u_ppwm/u_ex/state_q[2] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_tiehi \u_ppwm/u_ex/_1112__27  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net27));
 sg13g2_tiehi \u_ppwm/u_ex/_1122__28  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net28));
 sg13g2_tiehi \u_ppwm/u_ex/_1111__29  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net29));
 sg13g2_tiehi \u_ppwm/u_ex/_1118__30  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net30));
 sg13g2_tiehi \u_ppwm/u_ex/_1110__31  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net31));
 sg13g2_tiehi \u_ppwm/u_ex/_1126__32  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net32));
 sg13g2_tiehi \u_ppwm/u_ex/_1109__33  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_tiehi \u_ppwm/u_ex/_1117__34  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net34));
 sg13g2_tiehi \u_ppwm/u_ex/_1108__35  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net35));
 sg13g2_tiehi \u_ppwm/u_ex/_1121__36  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net36));
 sg13g2_tiehi \u_ppwm/u_ex/_1107__37  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_tiehi \u_ppwm/u_ex/_1116__38  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi \u_ppwm/u_ex/_1106__39  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi \u_ppwm/u_ex/_1123__40  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_tiehi \u_ppwm/u_ex/_1105__41  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net41));
 sg13g2_tiehi \u_ppwm/u_ex/_1115__42  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_tiehi \u_ppwm/u_ex/_1104__43  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_tiehi \u_ppwm/u_ex/_1120__44  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net44));
 sg13g2_tiehi \u_ppwm/u_ex/_1103__45  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net45));
 sg13g2_tiehi \u_ppwm/u_ex/_1114__46  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net46));
 sg13g2_tiehi \u_ppwm/u_ex/_1102__47  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net47));
 sg13g2_tiehi \u_ppwm/u_ex/_1127__48  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net48));
 sg13g2_tiehi \u_ppwm/u_ex/_1101__49  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net49));
 sg13g2_tiehi \u_ppwm/u_ex/_1113__50  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net50));
 sg13g2_tiehi \u_ppwm/u_ex/_1100__51  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net51));
 sg13g2_tiehi \u_ppwm/u_ex/_1099__52  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net52));
 sg13g2_tiehi \u_ppwm/u_ex/_1124__53  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net53));
 sg13g2_tiehi \u_ppwm/u_ex/_1125__54  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net54));
 sg13g2_tiehi \u_ppwm/u_mem/_1190__55  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net55));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_053_  (.VDD(VPWR),
    .Y(\u_ppwm/u_global_counter/_020_ ),
    .A(net599),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_054_  (.VDD(VPWR),
    .Y(\u_ppwm/u_global_counter/_021_ ),
    .A(\u_ppwm/global_counter[11] ),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_055_  (.VDD(VPWR),
    .Y(\u_ppwm/u_global_counter/_022_ ),
    .A(\u_ppwm/global_counter[13] ),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_056_  (.VDD(VPWR),
    .Y(\u_ppwm/u_global_counter/_023_ ),
    .A(net622),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_057_  (.VDD(VPWR),
    .Y(\u_ppwm/u_global_counter/_024_ ),
    .A(net645),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_058_  (.VDD(VPWR),
    .Y(\u_ppwm/u_global_counter/_025_ ),
    .A(net620),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_059_  (.VDD(VPWR),
    .Y(\u_ppwm/u_global_counter/_026_ ),
    .A(net398),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_060_  (.B(net398),
    .A(net445),
    .X(\u_ppwm/u_global_counter/_000_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_061_  (.B(net444),
    .C(net398),
    .A(net445),
    .Y(\u_ppwm/u_global_counter/_027_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_global_counter/_062_  (.A2(net399),
    .A1(net445),
    .B1(net444),
    .X(\u_ppwm/u_global_counter/_028_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_global_counter/_063_  (.A(\u_ppwm/u_global_counter/_027_ ),
    .B(\u_ppwm/u_global_counter/_028_ ),
    .X(\u_ppwm/u_global_counter/_001_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_064_  (.B(\u_ppwm/global_counter[1] ),
    .C(net443),
    .A(net445),
    .Y(\u_ppwm/u_global_counter/_029_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net398));
 sg13g2_xnor2_1 \u_ppwm/u_global_counter/_065_  (.Y(\u_ppwm/u_global_counter/_002_ ),
    .A(net443),
    .B(\u_ppwm/u_global_counter/_027_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_global_counter/_066_  (.A(\u_ppwm/u_global_counter/_020_ ),
    .B(\u_ppwm/u_global_counter/_029_ ),
    .Y(\u_ppwm/u_global_counter/_030_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_global_counter/_067_  (.Y(\u_ppwm/u_global_counter/_003_ ),
    .A(net599),
    .B(\u_ppwm/u_global_counter/_029_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_068_  (.B(\u_ppwm/u_global_counter/_030_ ),
    .A(net590),
    .X(\u_ppwm/u_global_counter/_004_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_069_  (.B(net599),
    .C(net590),
    .A(net659),
    .Y(\u_ppwm/u_global_counter/_031_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net627));
 sg13g2_nor2_1 \u_ppwm/u_global_counter/_070_  (.A(\u_ppwm/u_global_counter/_027_ ),
    .B(\u_ppwm/u_global_counter/_031_ ),
    .Y(\u_ppwm/u_global_counter/_032_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_071_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net590),
    .A2(\u_ppwm/u_global_counter/_030_ ),
    .Y(\u_ppwm/u_global_counter/_033_ ),
    .B1(net627));
 sg13g2_nor2_1 \u_ppwm/u_global_counter/_072_  (.A(\u_ppwm/u_global_counter/_032_ ),
    .B(net628),
    .Y(\u_ppwm/u_global_counter/_005_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_073_  (.B(\u_ppwm/u_global_counter/_032_ ),
    .A(net604),
    .X(\u_ppwm/u_global_counter/_006_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_074_  (.B(\u_ppwm/global_counter[1] ),
    .C(net604),
    .A(net653),
    .Y(\u_ppwm/u_global_counter/_034_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net630));
 sg13g2_nor3_2 \u_ppwm/u_global_counter/_075_  (.A(\u_ppwm/u_global_counter/_026_ ),
    .B(\u_ppwm/u_global_counter/_031_ ),
    .C(net666),
    .Y(\u_ppwm/u_global_counter/_035_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_076_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net604),
    .A2(\u_ppwm/u_global_counter/_032_ ),
    .Y(\u_ppwm/u_global_counter/_036_ ),
    .B1(net630));
 sg13g2_nor2_1 \u_ppwm/u_global_counter/_077_  (.A(\u_ppwm/u_global_counter/_035_ ),
    .B(net631),
    .Y(\u_ppwm/u_global_counter/_007_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_078_  (.B(\u_ppwm/u_global_counter/_035_ ),
    .A(net201),
    .X(\u_ppwm/u_global_counter/_008_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_079_  (.B(net441),
    .C(\u_ppwm/u_global_counter/_035_ ),
    .A(net442),
    .Y(\u_ppwm/u_global_counter/_037_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_global_counter/_080_  (.A2(\u_ppwm/u_global_counter/_035_ ),
    .A1(net201),
    .B1(net441),
    .X(\u_ppwm/u_global_counter/_038_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_global_counter/_081_  (.A(\u_ppwm/u_global_counter/_037_ ),
    .B(\u_ppwm/u_global_counter/_038_ ),
    .X(\u_ppwm/u_global_counter/_009_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_082_  (.B(net639),
    .C(net575),
    .A(net201),
    .Y(\u_ppwm/u_global_counter/_039_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_global_counter/_035_ ));
 sg13g2_xnor2_1 \u_ppwm/u_global_counter/_083_  (.Y(\u_ppwm/u_global_counter/_010_ ),
    .A(net575),
    .B(\u_ppwm/u_global_counter/_037_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_084_  (.B(net639),
    .C(net575),
    .A(net442),
    .Y(\u_ppwm/u_global_counter/_040_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/global_counter[11] ));
 sg13g2_nor3_1 \u_ppwm/u_global_counter/_085_  (.A(\u_ppwm/u_global_counter/_031_ ),
    .B(\u_ppwm/u_global_counter/_034_ ),
    .C(\u_ppwm/u_global_counter/_040_ ),
    .Y(\u_ppwm/u_global_counter/_041_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_global_counter/_086_  (.Y(\u_ppwm/u_global_counter/_011_ ),
    .B1(\u_ppwm/u_global_counter/_041_ ),
    .B2(net398),
    .A2(net640),
    .A1(\u_ppwm/u_global_counter/_021_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_087_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net398),
    .A2(net392),
    .Y(\u_ppwm/u_global_counter/_042_ ),
    .B1(net440));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_088_  (.B(net398),
    .C(net392),
    .A(net633),
    .Y(\u_ppwm/u_global_counter/_043_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_global_counter/_089_  (.A(\u_ppwm/u_global_counter/_042_ ),
    .B_N(\u_ppwm/u_global_counter/_043_ ),
    .Y(\u_ppwm/u_global_counter/_012_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 \u_ppwm/u_global_counter/_090_  (.X(\u_ppwm/u_global_counter/_044_ ),
    .A(net633),
    .B(\u_ppwm/global_counter[13] ),
    .C(net398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_global_counter/_091_  (.Y(\u_ppwm/u_global_counter/_013_ ),
    .B1(\u_ppwm/u_global_counter/_044_ ),
    .B2(net392),
    .A2(net634),
    .A1(\u_ppwm/u_global_counter/_022_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_092_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net392),
    .A2(\u_ppwm/u_global_counter/_044_ ),
    .Y(\u_ppwm/u_global_counter/_045_ ),
    .B1(net608));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_093_  (.B(\u_ppwm/u_global_counter/_041_ ),
    .C(\u_ppwm/u_global_counter/_044_ ),
    .A(net608),
    .Y(\u_ppwm/u_global_counter/_046_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_global_counter/_094_  (.A(net609),
    .B_N(\u_ppwm/u_global_counter/_046_ ),
    .Y(\u_ppwm/u_global_counter/_014_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 \u_ppwm/u_global_counter/_095_  (.X(\u_ppwm/u_global_counter/_047_ ),
    .A(net608),
    .B(net622),
    .C(\u_ppwm/u_global_counter/_044_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_global_counter/_096_  (.A(net392),
    .B(\u_ppwm/u_global_counter/_047_ ),
    .X(\u_ppwm/u_global_counter/_048_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_097_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_global_counter/_023_ ),
    .A2(\u_ppwm/u_global_counter/_046_ ),
    .Y(\u_ppwm/u_global_counter/_015_ ),
    .B1(\u_ppwm/u_global_counter/_048_ ));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_098_  (.B(net392),
    .C(\u_ppwm/u_global_counter/_047_ ),
    .A(net439),
    .Y(\u_ppwm/u_global_counter/_049_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_099_  (.B(\u_ppwm/u_global_counter/_048_ ),
    .A(net439),
    .X(\u_ppwm/u_global_counter/_016_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_global_counter/_100_  (.A(net439),
    .B(net645),
    .X(\u_ppwm/u_global_counter/_050_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_101_  (.B(\u_ppwm/u_global_counter/_047_ ),
    .C(\u_ppwm/u_global_counter/_050_ ),
    .A(net392),
    .Y(\u_ppwm/u_global_counter/_051_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 \u_ppwm/u_global_counter/_102_  (.Y(\u_ppwm/u_global_counter/_017_ ),
    .B1(\u_ppwm/u_global_counter/_050_ ),
    .B2(\u_ppwm/u_global_counter/_048_ ),
    .A2(\u_ppwm/u_global_counter/_049_ ),
    .A1(\u_ppwm/u_global_counter/_024_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 \u_ppwm/u_global_counter/_103_  (.A(net620),
    .B(net392),
    .C(\u_ppwm/u_global_counter/_047_ ),
    .D(\u_ppwm/u_global_counter/_050_ ),
    .X(\u_ppwm/u_global_counter/_052_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_104_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_global_counter/_025_ ),
    .A2(\u_ppwm/u_global_counter/_051_ ),
    .Y(\u_ppwm/u_global_counter/_018_ ),
    .B1(\u_ppwm/u_global_counter/_052_ ));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_105_  (.B(\u_ppwm/u_global_counter/_052_ ),
    .A(net585),
    .X(\u_ppwm/u_global_counter/_019_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_106_  (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_global_counter/_000_ ),
    .Q(\u_ppwm/global_counter[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_107_  (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_global_counter/_001_ ),
    .Q(\u_ppwm/global_counter[1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_global_counter/_108_  (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net656),
    .Q(\u_ppwm/global_counter[2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_109_  (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net600),
    .Q(\u_ppwm/global_counter[3] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_110_  (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net591),
    .Q(\u_ppwm/global_counter[4] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_111_  (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net629),
    .Q(\u_ppwm/global_counter[5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_112_  (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net605),
    .Q(\u_ppwm/global_counter[6] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_113_  (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net632),
    .Q(\u_ppwm/global_counter[7] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_114_  (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net202),
    .Q(\u_ppwm/global_counter[8] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_115_  (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_global_counter/_009_ ),
    .Q(\u_ppwm/global_counter[9] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_116_  (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net576),
    .Q(\u_ppwm/global_counter[10] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_117_  (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net641),
    .Q(\u_ppwm/global_counter[11] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_118_  (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_global_counter/_012_ ),
    .Q(\u_ppwm/global_counter[12] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_119_  (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net635),
    .Q(\u_ppwm/global_counter[13] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_120_  (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net610),
    .Q(\u_ppwm/global_counter[14] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_121_  (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net623),
    .Q(\u_ppwm/global_counter[15] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_122_  (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_global_counter/_016_ ),
    .Q(\u_ppwm/global_counter[16] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_123_  (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net646),
    .Q(\u_ppwm/global_counter[17] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_124_  (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net621),
    .Q(\u_ppwm/global_counter[18] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_125_  (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net586),
    .Q(\u_ppwm/global_counter[19] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_inv_1 \u_ppwm/u_mem/_0613_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0126_ ),
    .A(net535),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0614_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0127_ ),
    .A(net1),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0615_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0128_ ),
    .A(net295),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0616_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0129_ ),
    .A(net527),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0617_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0130_ ),
    .A(net222),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0618_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0131_ ),
    .A(net290),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0619_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0132_ ),
    .A(net307),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0620_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0133_ ),
    .A(net343),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0621_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0134_ ),
    .A(net537),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0622_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0135_ ),
    .A(net528),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0623_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0136_ ),
    .A(net318),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0624_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0137_ ),
    .A(net253),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0625_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0138_ ),
    .A(net258),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0626_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0139_ ),
    .A(net301),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0627_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0140_ ),
    .A(net312),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0628_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0141_ ),
    .A(net328),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0629_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0142_ ),
    .A(net213),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0630_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0143_ ),
    .A(net339),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0631_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0144_ ),
    .A(net520),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0632_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0145_ ),
    .A(net582),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0633_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0146_ ),
    .A(net526),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0634_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0147_ ),
    .A(net205),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0635_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0148_ ),
    .A(net257),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0636_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0149_ ),
    .A(net232),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0637_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0150_ ),
    .A(net305),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0638_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0151_ ),
    .A(net230),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0639_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0152_ ),
    .A(net568),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0640_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0153_ ),
    .A(net538),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0641_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0154_ ),
    .A(net571),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0642_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0155_ ),
    .A(net326),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0643_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0156_ ),
    .A(net580),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0644_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0157_ ),
    .A(net319),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0645_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0158_ ),
    .A(net236),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0646_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0159_ ),
    .A(net249),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0647_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0160_ ),
    .A(net322),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0648_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0161_ ),
    .A(net583),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0649_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0162_ ),
    .A(net345),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0650_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0163_ ),
    .A(net540),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0651_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0164_ ),
    .A(net244),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0652_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0165_ ),
    .A(net234),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0653_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0166_ ),
    .A(net255),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0654_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0167_ ),
    .A(net265),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0655_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0168_ ),
    .A(net348),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0656_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0169_ ),
    .A(net579),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0657_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0170_ ),
    .A(net297),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0658_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0171_ ),
    .A(net292),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0659_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0172_ ),
    .A(net228),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0660_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0173_ ),
    .A(net303),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0661_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0174_ ),
    .A(net251),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0662_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0175_ ),
    .A(net267),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0663_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0176_ ),
    .A(net592),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0664_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0177_ ),
    .A(net306),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0665_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0178_ ),
    .A(net264),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0666_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0179_ ),
    .A(net224),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0667_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0180_ ),
    .A(net315),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0668_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0181_ ),
    .A(net531),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0669_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0182_ ),
    .A(net286),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0670_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0183_ ),
    .A(net317),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0671_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0184_ ),
    .A(net271),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0672_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0185_ ),
    .A(net553),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0673_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0186_ ),
    .A(net536),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0674_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0187_ ),
    .A(net245),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0675_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0188_ ),
    .A(net541),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0676_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0189_ ),
    .A(net309),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0677_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0190_ ),
    .A(net240),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0678_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0191_ ),
    .A(net269),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0679_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0192_ ),
    .A(net542),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0680_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0193_ ),
    .A(net278),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0681_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0194_ ),
    .A(net310),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0682_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0195_ ),
    .A(net522),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0683_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0196_ ),
    .A(net556),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0684_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0197_ ),
    .A(net596),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0685_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0198_ ),
    .A(net273),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0686_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0199_ ),
    .A(net335),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0687_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0200_ ),
    .A(net320),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0688_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0201_ ),
    .A(net337),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0689_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0202_ ),
    .A(net220),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0690_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0203_ ),
    .A(net545),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0691_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0204_ ),
    .A(net314),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0692_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0205_ ),
    .A(net226),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0693_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0206_ ),
    .A(net559),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0694_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0207_ ),
    .A(net324),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0695_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0208_ ),
    .A(net554),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0696_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0209_ ),
    .A(net329),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0697_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0210_ ),
    .A(net288),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0698_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0211_ ),
    .A(net570),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0699_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0212_ ),
    .A(net336),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0700_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0213_ ),
    .A(net262),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0701_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0214_ ),
    .A(net581),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0702_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0215_ ),
    .A(net524),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0703_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0216_ ),
    .A(net282),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0704_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0217_ ),
    .A(net347),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0705_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0218_ ),
    .A(net331),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0706_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0219_ ),
    .A(net529),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0707_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0220_ ),
    .A(net558),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0708_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0221_ ),
    .A(net543),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0709_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0222_ ),
    .A(net551),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0710_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0223_ ),
    .A(net564),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0711_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0224_ ),
    .A(net275),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0712_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0225_ ),
    .A(net293),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0713_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0226_ ),
    .A(net532),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0714_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0227_ ),
    .A(net280),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0715_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0228_ ),
    .A(net563),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0716_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0229_ ),
    .A(net561),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0717_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0230_ ),
    .A(net298),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0718_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0231_ ),
    .A(net284),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0719_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0232_ ),
    .A(net560),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0720_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0233_ ),
    .A(net277),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0721_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0234_ ),
    .A(net242),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0722_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0235_ ),
    .A(net341),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0723_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0236_ ),
    .A(net577),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0724_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0237_ ),
    .A(\u_ppwm/u_mem/memory[1] ),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_mem/_0725_  (.Y(\u_ppwm/u_mem/_0238_ ),
    .A(net488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0726_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0239_ ),
    .A(net333),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0727_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0240_ ),
    .A(net475),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_mem/_0728_  (.VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0241_ ),
    .A(\u_ppwm/pc[2] ),
    .VSS(VGND));
 sg13g2_inv_4 \u_ppwm/u_mem/_0729_  (.A(net467),
    .Y(\u_ppwm/u_mem/_0242_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_mem/_0730_  (.A(\u_ppwm/u_mem/_0127_ ),
    .B(\u_ppwm/u_mem/_0238_ ),
    .C(\u_ppwm/mem_write_done ),
    .Y(\u_ppwm/u_mem/_0243_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_mem/_0731_  (.A(net1),
    .B(\u_ppwm/u_mem/_0238_ ),
    .Y(\u_ppwm/u_mem/_0244_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0732_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0239_ ),
    .A2(\u_ppwm/u_mem/_0244_ ),
    .Y(\u_ppwm/u_mem/_0004_ ),
    .B1(\u_ppwm/u_mem/_0243_ ));
 sg13g2_nand3_1 \u_ppwm/u_mem/_0733_  (.B(net587),
    .C(net606),
    .A(net565),
    .Y(\u_ppwm/u_mem/_0245_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_mem/_0734_  (.B(\u_ppwm/u_mem/bit_count[1] ),
    .C(net617),
    .A(net611),
    .Y(\u_ppwm/u_mem/_0246_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_mem/_0735_  (.A(net618),
    .B(\u_ppwm/u_mem/_0245_ ),
    .C(\u_ppwm/u_mem/_0246_ ),
    .Y(\u_ppwm/u_mem/_0247_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0736_  (.Y(\u_ppwm/u_mem/_0248_ ),
    .A(net400),
    .B(net488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 \u_ppwm/u_mem/_0737_  (.A(net618),
    .B(\u_ppwm/u_mem/_0245_ ),
    .C(\u_ppwm/u_mem/_0246_ ),
    .D(\u_ppwm/u_mem/_0248_ ),
    .Y(\u_ppwm/u_mem/_0249_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 \u_ppwm/u_mem/_0738_  (.A2(\u_ppwm/u_mem/_0244_ ),
    .A1(net625),
    .B1(\u_ppwm/u_mem/_0249_ ),
    .X(\u_ppwm/u_mem/_0005_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_mem/_0739_  (.B(net488),
    .C(net333),
    .A(net1),
    .Y(\u_ppwm/u_mem/_0250_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0740_  (.B1(\u_ppwm/u_mem/_0250_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0006_ ),
    .VSS(VGND),
    .A1(net619),
    .A2(\u_ppwm/u_mem/_0248_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0741_  (.A0(\u_ppwm/u_mem/memory[70] ),
    .A1(\u_ppwm/u_mem/memory[77] ),
    .S(net478),
    .X(\u_ppwm/u_mem/_0251_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0742_  (.A0(\u_ppwm/u_mem/memory[56] ),
    .A1(\u_ppwm/u_mem/memory[63] ),
    .S(net481),
    .X(\u_ppwm/u_mem/_0252_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0743_  (.Y(\u_ppwm/u_mem/_0253_ ),
    .A(net396),
    .B(\u_ppwm/u_mem/_0252_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0744_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net472),
    .A2(\u_ppwm/u_mem/_0251_ ),
    .Y(\u_ppwm/u_mem/_0254_ ),
    .B1(net470));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0745_  (.A0(\u_ppwm/u_mem/memory[84] ),
    .A1(\u_ppwm/u_mem/memory[91] ),
    .S(net477),
    .X(\u_ppwm/u_mem/_0255_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0746_  (.Y(\u_ppwm/u_mem/_0256_ ),
    .A(net395),
    .B(\u_ppwm/u_mem/_0255_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0747_  (.A0(\u_ppwm/u_mem/memory[98] ),
    .A1(\u_ppwm/u_mem/memory[105] ),
    .S(net477),
    .X(\u_ppwm/u_mem/_0257_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0748_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net472),
    .A2(\u_ppwm/u_mem/_0257_ ),
    .Y(\u_ppwm/u_mem/_0258_ ),
    .B1(net394));
 sg13g2_a221oi_1 \u_ppwm/u_mem/_0749_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_mem/_0258_ ),
    .C1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0256_ ),
    .A1(\u_ppwm/u_mem/_0253_ ),
    .Y(\u_ppwm/u_mem/_0259_ ),
    .A2(\u_ppwm/u_mem/_0254_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0750_  (.S0(net484),
    .A0(\u_ppwm/u_mem/memory[0] ),
    .A1(\u_ppwm/u_mem/memory[7] ),
    .A2(\u_ppwm/u_mem/memory[14] ),
    .A3(\u_ppwm/u_mem/memory[21] ),
    .S1(net475),
    .X(\u_ppwm/u_mem/_0260_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_mem/_0751_  (.Y(\u_ppwm/u_mem/_0261_ ),
    .B(\u_ppwm/u_mem/_0241_ ),
    .A_N(\u_ppwm/u_mem/_0260_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0752_  (.A0(\u_ppwm/u_mem/memory[42] ),
    .A1(\u_ppwm/u_mem/memory[49] ),
    .S(net486),
    .X(\u_ppwm/u_mem/_0262_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0753_  (.A0(\u_ppwm/u_mem/memory[28] ),
    .A1(\u_ppwm/u_mem/memory[35] ),
    .S(net483),
    .X(\u_ppwm/u_mem/_0263_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0754_  (.Y(\u_ppwm/u_mem/_0264_ ),
    .A(net397),
    .B(\u_ppwm/u_mem/_0263_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0755_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net473),
    .A2(\u_ppwm/u_mem/_0262_ ),
    .Y(\u_ppwm/u_mem/_0265_ ),
    .B1(net393));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0756_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0264_ ),
    .A2(\u_ppwm/u_mem/_0265_ ),
    .Y(\u_ppwm/u_mem/_0266_ ),
    .B1(net467));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0757_  (.A2(\u_ppwm/u_mem/_0266_ ),
    .A1(\u_ppwm/u_mem/_0261_ ),
    .B1(\u_ppwm/u_mem/_0259_ ),
    .X(\u_ppwm/instr[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0758_  (.A0(\u_ppwm/u_mem/memory[99] ),
    .A1(\u_ppwm/u_mem/memory[106] ),
    .S(net477),
    .X(\u_ppwm/u_mem/_0267_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0759_  (.A0(\u_ppwm/u_mem/memory[85] ),
    .A1(\u_ppwm/u_mem/memory[92] ),
    .S(net477),
    .X(\u_ppwm/u_mem/_0268_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0760_  (.Y(\u_ppwm/u_mem/_0269_ ),
    .A(net395),
    .B(\u_ppwm/u_mem/_0268_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0761_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net472),
    .A2(\u_ppwm/u_mem/_0267_ ),
    .Y(\u_ppwm/u_mem/_0270_ ),
    .B1(net394));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0762_  (.S0(net478),
    .A0(\u_ppwm/u_mem/memory[57] ),
    .A1(\u_ppwm/u_mem/memory[64] ),
    .A2(\u_ppwm/u_mem/memory[71] ),
    .A3(\u_ppwm/u_mem/memory[78] ),
    .S1(net472),
    .X(\u_ppwm/u_mem/_0271_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0763_  (.B1(net467),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0272_ ),
    .VSS(VGND),
    .A1(net470),
    .A2(\u_ppwm/u_mem/_0271_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0764_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0269_ ),
    .A2(\u_ppwm/u_mem/_0270_ ),
    .Y(\u_ppwm/u_mem/_0273_ ),
    .B1(\u_ppwm/u_mem/_0272_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0765_  (.Y(\u_ppwm/u_mem/_0274_ ),
    .A(\u_ppwm/u_mem/memory[36] ),
    .B(net483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0766_  (.B1(\u_ppwm/u_mem/_0274_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0275_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0209_ ),
    .A2(net483));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0767_  (.Y(\u_ppwm/u_mem/_0276_ ),
    .A(\u_ppwm/u_mem/memory[50] ),
    .B(net482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0768_  (.B1(\u_ppwm/u_mem/_0276_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0277_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0195_ ),
    .A2(net482));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0769_  (.Y(\u_ppwm/u_mem/_0278_ ),
    .A(\u_ppwm/u_mem/memory[22] ),
    .B(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0770_  (.B1(\u_ppwm/u_mem/_0278_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0279_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0223_ ),
    .A2(net484));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0771_  (.Y(\u_ppwm/u_mem/_0280_ ),
    .A(\u_ppwm/u_mem/memory[8] ),
    .B(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0772_  (.B1(\u_ppwm/u_mem/_0280_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0281_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0237_ ),
    .A2(net484));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0773_  (.S0(net475),
    .A0(\u_ppwm/u_mem/_0275_ ),
    .A1(\u_ppwm/u_mem/_0277_ ),
    .A2(\u_ppwm/u_mem/_0281_ ),
    .A3(\u_ppwm/u_mem/_0279_ ),
    .S1(net393),
    .X(\u_ppwm/u_mem/_0282_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0774_  (.A2(\u_ppwm/u_mem/_0282_ ),
    .A1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0273_ ),
    .X(\u_ppwm/instr[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0775_  (.A0(\u_ppwm/u_mem/memory[100] ),
    .A1(\u_ppwm/u_mem/memory[107] ),
    .S(net477),
    .X(\u_ppwm/u_mem/_0283_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0776_  (.Y(\u_ppwm/u_mem/_0284_ ),
    .A(net471),
    .B(\u_ppwm/u_mem/_0283_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0777_  (.A0(\u_ppwm/u_mem/memory[86] ),
    .A1(\u_ppwm/u_mem/memory[93] ),
    .S(net480),
    .X(\u_ppwm/u_mem/_0285_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0778_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net395),
    .A2(\u_ppwm/u_mem/_0285_ ),
    .Y(\u_ppwm/u_mem/_0286_ ),
    .B1(net394));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0779_  (.A0(\u_ppwm/u_mem/memory[72] ),
    .A1(\u_ppwm/u_mem/memory[79] ),
    .S(net478),
    .X(\u_ppwm/u_mem/_0287_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0780_  (.Y(\u_ppwm/u_mem/_0288_ ),
    .A(net471),
    .B(\u_ppwm/u_mem/_0287_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0781_  (.A0(\u_ppwm/u_mem/memory[58] ),
    .A1(\u_ppwm/u_mem/memory[65] ),
    .S(net478),
    .X(\u_ppwm/u_mem/_0289_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0782_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net395),
    .A2(\u_ppwm/u_mem/_0289_ ),
    .Y(\u_ppwm/u_mem/_0290_ ),
    .B1(net470));
 sg13g2_a221oi_1 \u_ppwm/u_mem/_0783_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_mem/_0290_ ),
    .C1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0288_ ),
    .A1(\u_ppwm/u_mem/_0284_ ),
    .Y(\u_ppwm/u_mem/_0291_ ),
    .A2(\u_ppwm/u_mem/_0286_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0784_  (.Y(\u_ppwm/u_mem/_0292_ ),
    .A(\u_ppwm/u_mem/memory[37] ),
    .B(net486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0785_  (.B1(\u_ppwm/u_mem/_0292_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0293_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0208_ ),
    .A2(net486));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0786_  (.Y(\u_ppwm/u_mem/_0294_ ),
    .A(\u_ppwm/u_mem/memory[51] ),
    .B(net482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0787_  (.B1(\u_ppwm/u_mem/_0294_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0295_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0194_ ),
    .A2(net482));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0788_  (.Y(\u_ppwm/u_mem/_0296_ ),
    .A(\u_ppwm/u_mem/memory[23] ),
    .B(net485),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0789_  (.B1(\u_ppwm/u_mem/_0296_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0297_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0222_ ),
    .A2(net485));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0790_  (.Y(\u_ppwm/u_mem/_0298_ ),
    .A(\u_ppwm/u_mem/memory[9] ),
    .B(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0791_  (.B1(\u_ppwm/u_mem/_0298_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0299_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0236_ ),
    .A2(net484));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0792_  (.S0(net475),
    .A0(\u_ppwm/u_mem/_0293_ ),
    .A1(\u_ppwm/u_mem/_0295_ ),
    .A2(\u_ppwm/u_mem/_0299_ ),
    .A3(\u_ppwm/u_mem/_0297_ ),
    .S1(net393),
    .X(\u_ppwm/u_mem/_0300_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0793_  (.A2(\u_ppwm/u_mem/_0300_ ),
    .A1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0291_ ),
    .X(\u_ppwm/instr[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0794_  (.A0(\u_ppwm/u_mem/memory[101] ),
    .A1(\u_ppwm/u_mem/_0000_ ),
    .S(net476),
    .X(\u_ppwm/u_mem/_0301_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0795_  (.Y(\u_ppwm/u_mem/_0302_ ),
    .A(net471),
    .B(\u_ppwm/u_mem/_0301_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0796_  (.A0(\u_ppwm/u_mem/memory[87] ),
    .A1(\u_ppwm/u_mem/memory[94] ),
    .S(net480),
    .X(\u_ppwm/u_mem/_0303_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0797_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net395),
    .A2(\u_ppwm/u_mem/_0303_ ),
    .Y(\u_ppwm/u_mem/_0304_ ),
    .B1(net394));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0798_  (.A0(\u_ppwm/u_mem/memory[73] ),
    .A1(\u_ppwm/u_mem/memory[80] ),
    .S(net478),
    .X(\u_ppwm/u_mem/_0305_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0799_  (.Y(\u_ppwm/u_mem/_0306_ ),
    .A(net472),
    .B(\u_ppwm/u_mem/_0305_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0800_  (.A0(\u_ppwm/u_mem/memory[59] ),
    .A1(\u_ppwm/u_mem/memory[66] ),
    .S(net478),
    .X(\u_ppwm/u_mem/_0307_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0801_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net395),
    .A2(\u_ppwm/u_mem/_0307_ ),
    .Y(\u_ppwm/u_mem/_0308_ ),
    .B1(net470));
 sg13g2_a221oi_1 \u_ppwm/u_mem/_0802_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_mem/_0308_ ),
    .C1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0306_ ),
    .A1(\u_ppwm/u_mem/_0302_ ),
    .Y(\u_ppwm/u_mem/_0309_ ),
    .A2(\u_ppwm/u_mem/_0304_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0803_  (.A0(\u_ppwm/u_mem/_0207_ ),
    .A1(\u_ppwm/u_mem/_0200_ ),
    .S(net482),
    .X(\u_ppwm/u_mem/_0310_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0804_  (.A0(\u_ppwm/u_mem/memory[45] ),
    .A1(\u_ppwm/u_mem/memory[52] ),
    .S(net482),
    .X(\u_ppwm/u_mem/_0311_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0805_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net473),
    .A2(\u_ppwm/u_mem/_0311_ ),
    .Y(\u_ppwm/u_mem/_0312_ ),
    .B1(net393));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0806_  (.B1(\u_ppwm/u_mem/_0312_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0313_ ),
    .VSS(VGND),
    .A1(net473),
    .A2(\u_ppwm/u_mem/_0310_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0807_  (.S0(net397),
    .A0(\u_ppwm/u_mem/_0221_ ),
    .A1(\u_ppwm/u_mem/_0235_ ),
    .A2(\u_ppwm/u_mem/_0214_ ),
    .A3(\u_ppwm/u_mem/_0228_ ),
    .S1(net485),
    .X(\u_ppwm/u_mem/_0314_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0808_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net393),
    .A2(\u_ppwm/u_mem/_0314_ ),
    .Y(\u_ppwm/u_mem/_0315_ ),
    .B1(net467));
 sg13g2_a21o_1 \u_ppwm/u_mem/_0809_  (.A2(\u_ppwm/u_mem/_0315_ ),
    .A1(\u_ppwm/u_mem/_0313_ ),
    .B1(\u_ppwm/u_mem/_0309_ ),
    .X(\u_ppwm/instr[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0810_  (.B1(net471),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0316_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/memory[102] ),
    .A2(net476));
 sg13g2_a21o_1 \u_ppwm/u_mem/_0811_  (.A2(net476),
    .A1(\u_ppwm/u_mem/_0129_ ),
    .B1(\u_ppwm/u_mem/_0316_ ),
    .X(\u_ppwm/u_mem/_0317_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0812_  (.A0(\u_ppwm/u_mem/memory[88] ),
    .A1(\u_ppwm/u_mem/memory[95] ),
    .S(net480),
    .X(\u_ppwm/u_mem/_0318_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0813_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net396),
    .A2(\u_ppwm/u_mem/_0318_ ),
    .Y(\u_ppwm/u_mem/_0319_ ),
    .B1(net394));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0814_  (.S0(net478),
    .A0(\u_ppwm/u_mem/memory[60] ),
    .A1(\u_ppwm/u_mem/memory[67] ),
    .A2(\u_ppwm/u_mem/memory[74] ),
    .A3(\u_ppwm/u_mem/memory[81] ),
    .S1(net472),
    .X(\u_ppwm/u_mem/_0320_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0815_  (.B1(net467),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0321_ ),
    .VSS(VGND),
    .A1(net470),
    .A2(\u_ppwm/u_mem/_0320_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0816_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0317_ ),
    .A2(\u_ppwm/u_mem/_0319_ ),
    .Y(\u_ppwm/u_mem/_0322_ ),
    .B1(\u_ppwm/u_mem/_0321_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0817_  (.A0(\u_ppwm/u_mem/memory[18] ),
    .A1(\u_ppwm/u_mem/memory[25] ),
    .S(net485),
    .X(\u_ppwm/u_mem/_0323_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0818_  (.Y(\u_ppwm/u_mem/_0324_ ),
    .A(net475),
    .B(\u_ppwm/u_mem/_0323_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0819_  (.A0(\u_ppwm/u_mem/memory[4] ),
    .A1(\u_ppwm/u_mem/memory[11] ),
    .S(net485),
    .X(\u_ppwm/u_mem/_0325_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0820_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net397),
    .A2(\u_ppwm/u_mem/_0325_ ),
    .Y(\u_ppwm/u_mem/_0326_ ),
    .B1(net469));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0821_  (.B1(net474),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0327_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/memory[46] ),
    .A2(net482));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0822_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0185_ ),
    .A2(net482),
    .Y(\u_ppwm/u_mem/_0328_ ),
    .B1(\u_ppwm/u_mem/_0327_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0823_  (.A0(\u_ppwm/u_mem/memory[32] ),
    .A1(\u_ppwm/u_mem/memory[39] ),
    .S(net481),
    .X(\u_ppwm/u_mem/_0329_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0824_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net396),
    .A2(\u_ppwm/u_mem/_0329_ ),
    .Y(\u_ppwm/u_mem/_0330_ ),
    .B1(net393));
 sg13g2_nand2b_1 \u_ppwm/u_mem/_0825_  (.Y(\u_ppwm/u_mem/_0331_ ),
    .B(\u_ppwm/u_mem/_0330_ ),
    .A_N(\u_ppwm/u_mem/_0328_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0826_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0324_ ),
    .A2(\u_ppwm/u_mem/_0326_ ),
    .Y(\u_ppwm/u_mem/_0332_ ),
    .B1(net467));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0827_  (.A2(\u_ppwm/u_mem/_0332_ ),
    .A1(\u_ppwm/u_mem/_0331_ ),
    .B1(\u_ppwm/u_mem/_0322_ ),
    .X(\u_ppwm/instr[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_mem/_0828_  (.A(\u_ppwm/u_mem/_0002_ ),
    .B_N(net476),
    .Y(\u_ppwm/u_mem/_0333_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0829_  (.B1(net471),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0334_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/memory[103] ),
    .A2(net476));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0830_  (.Y(\u_ppwm/u_mem/_0335_ ),
    .A(\u_ppwm/u_mem/memory[96] ),
    .B(net480),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_mem/_0831_  (.Y(\u_ppwm/u_mem/_0336_ ),
    .B(\u_ppwm/u_mem/memory[89] ),
    .A_N(net480),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0832_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0335_ ),
    .A2(\u_ppwm/u_mem/_0336_ ),
    .Y(\u_ppwm/u_mem/_0337_ ),
    .B1(net472));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0833_  (.B1(net470),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0338_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0333_ ),
    .A2(\u_ppwm/u_mem/_0334_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0834_  (.S0(net478),
    .A0(\u_ppwm/u_mem/memory[61] ),
    .A1(\u_ppwm/u_mem/memory[68] ),
    .A2(\u_ppwm/u_mem/memory[75] ),
    .A3(\u_ppwm/u_mem/memory[82] ),
    .S1(net471),
    .X(\u_ppwm/u_mem/_0339_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_mem/_0835_  (.A(net470),
    .B(\u_ppwm/u_mem/_0339_ ),
    .Y(\u_ppwm/u_mem/_0340_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0836_  (.B1(net467),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0341_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0337_ ),
    .A2(\u_ppwm/u_mem/_0338_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0837_  (.A0(\u_ppwm/u_mem/memory[33] ),
    .A1(\u_ppwm/u_mem/memory[40] ),
    .S(net480),
    .X(\u_ppwm/u_mem/_0342_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0838_  (.A0(\u_ppwm/u_mem/memory[47] ),
    .A1(\u_ppwm/u_mem/memory[54] ),
    .S(net481),
    .X(\u_ppwm/u_mem/_0343_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0839_  (.A0(\u_ppwm/u_mem/memory[19] ),
    .A1(\u_ppwm/u_mem/memory[26] ),
    .S(net485),
    .X(\u_ppwm/u_mem/_0344_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0840_  (.A0(\u_ppwm/u_mem/memory[5] ),
    .A1(\u_ppwm/u_mem/memory[12] ),
    .S(net485),
    .X(\u_ppwm/u_mem/_0345_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0841_  (.S0(net474),
    .A0(\u_ppwm/u_mem/_0342_ ),
    .A1(\u_ppwm/u_mem/_0343_ ),
    .A2(\u_ppwm/u_mem/_0345_ ),
    .A3(\u_ppwm/u_mem/_0344_ ),
    .S1(net393),
    .X(\u_ppwm/u_mem/_0346_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0842_  (.Y(\u_ppwm/u_mem/_0347_ ),
    .A(\u_ppwm/u_mem/_0242_ ),
    .B(\u_ppwm/u_mem/_0346_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0843_  (.B1(\u_ppwm/u_mem/_0347_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/instr[5] ),
    .VSS(VGND),
    .A1(\u_ppwm/u_mem/_0340_ ),
    .A2(\u_ppwm/u_mem/_0341_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0844_  (.A0(\u_ppwm/u_mem/memory[76] ),
    .A1(\u_ppwm/u_mem/memory[83] ),
    .S(net476),
    .X(\u_ppwm/u_mem/_0348_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0845_  (.Y(\u_ppwm/u_mem/_0349_ ),
    .A(net471),
    .B(\u_ppwm/u_mem/_0348_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0846_  (.A0(\u_ppwm/u_mem/memory[62] ),
    .A1(\u_ppwm/u_mem/memory[69] ),
    .S(net479),
    .X(\u_ppwm/u_mem/_0350_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0847_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net395),
    .A2(\u_ppwm/u_mem/_0350_ ),
    .Y(\u_ppwm/u_mem/_0351_ ),
    .B1(net470));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0848_  (.A0(\u_ppwm/u_mem/memory[90] ),
    .A1(\u_ppwm/u_mem/memory[97] ),
    .S(net476),
    .X(\u_ppwm/u_mem/_0352_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0849_  (.A0(\u_ppwm/u_mem/memory[104] ),
    .A1(\u_ppwm/u_mem/_0003_ ),
    .S(net476),
    .X(\u_ppwm/u_mem/_0353_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0850_  (.Y(\u_ppwm/u_mem/_0354_ ),
    .A(net471),
    .B(\u_ppwm/u_mem/_0353_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0851_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net395),
    .A2(\u_ppwm/u_mem/_0352_ ),
    .Y(\u_ppwm/u_mem/_0355_ ),
    .B1(net394));
 sg13g2_a221oi_1 \u_ppwm/u_mem/_0852_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_mem/_0355_ ),
    .C1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0354_ ),
    .A1(\u_ppwm/u_mem/_0349_ ),
    .Y(\u_ppwm/u_mem/_0356_ ),
    .A2(\u_ppwm/u_mem/_0351_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0853_  (.A0(\u_ppwm/u_mem/_0204_ ),
    .A1(\u_ppwm/u_mem/_0197_ ),
    .S(net481),
    .X(\u_ppwm/u_mem/_0357_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0854_  (.A0(\u_ppwm/u_mem/memory[48] ),
    .A1(\u_ppwm/u_mem/memory[55] ),
    .S(net480),
    .X(\u_ppwm/u_mem/_0358_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0855_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net474),
    .A2(\u_ppwm/u_mem/_0358_ ),
    .Y(\u_ppwm/u_mem/_0359_ ),
    .B1(net394));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0856_  (.B1(\u_ppwm/u_mem/_0359_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0360_ ),
    .VSS(VGND),
    .A1(net474),
    .A2(\u_ppwm/u_mem/_0357_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0857_  (.S0(net397),
    .A0(\u_ppwm/u_mem/_0218_ ),
    .A1(\u_ppwm/u_mem/_0232_ ),
    .A2(\u_ppwm/u_mem/_0211_ ),
    .A3(\u_ppwm/u_mem/_0225_ ),
    .S1(net484),
    .X(\u_ppwm/u_mem/_0361_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0858_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net393),
    .A2(\u_ppwm/u_mem/_0361_ ),
    .Y(\u_ppwm/u_mem/_0362_ ),
    .B1(net467));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0859_  (.A2(\u_ppwm/u_mem/_0362_ ),
    .A1(\u_ppwm/u_mem/_0360_ ),
    .B1(\u_ppwm/u_mem/_0356_ ),
    .X(\u_ppwm/instr[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0860_  (.B1(net513),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0363_ ),
    .VSS(VGND),
    .A1(net423),
    .A2(net597));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0861_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net424),
    .A2(\u_ppwm/u_mem/_0237_ ),
    .Y(\u_ppwm/u_mem/_0007_ ),
    .B1(\u_ppwm/u_mem/_0363_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0862_  (.B1(net514),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0364_ ),
    .VSS(VGND),
    .A1(net434),
    .A2(\u_ppwm/u_mem/memory[1] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0863_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net434),
    .A2(\u_ppwm/u_mem/_0236_ ),
    .Y(\u_ppwm/u_mem/_0008_ ),
    .B1(\u_ppwm/u_mem/_0364_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0864_  (.B1(net516),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0365_ ),
    .VSS(VGND),
    .A1(net433),
    .A2(\u_ppwm/u_mem/memory[2] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0865_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net435),
    .A2(\u_ppwm/u_mem/_0235_ ),
    .Y(\u_ppwm/u_mem/_0009_ ),
    .B1(\u_ppwm/u_mem/_0365_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0866_  (.B1(net516),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0366_ ),
    .VSS(VGND),
    .A1(net437),
    .A2(\u_ppwm/u_mem/memory[3] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0867_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net437),
    .A2(\u_ppwm/u_mem/_0234_ ),
    .Y(\u_ppwm/u_mem/_0010_ ),
    .B1(\u_ppwm/u_mem/_0366_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0868_  (.B1(net515),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0367_ ),
    .VSS(VGND),
    .A1(net433),
    .A2(net242));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0869_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net433),
    .A2(\u_ppwm/u_mem/_0233_ ),
    .Y(\u_ppwm/u_mem/_0011_ ),
    .B1(\u_ppwm/u_mem/_0367_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0870_  (.B1(net515),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0368_ ),
    .VSS(VGND),
    .A1(net432),
    .A2(net277));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0871_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net432),
    .A2(\u_ppwm/u_mem/_0232_ ),
    .Y(\u_ppwm/u_mem/_0012_ ),
    .B1(\u_ppwm/u_mem/_0368_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0872_  (.B1(net513),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0369_ ),
    .VSS(VGND),
    .A1(net423),
    .A2(\u_ppwm/u_mem/memory[6] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0873_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net423),
    .A2(\u_ppwm/u_mem/_0231_ ),
    .Y(\u_ppwm/u_mem/_0013_ ),
    .B1(\u_ppwm/u_mem/_0369_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0874_  (.B1(net513),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0370_ ),
    .VSS(VGND),
    .A1(net423),
    .A2(net284));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0875_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net423),
    .A2(\u_ppwm/u_mem/_0230_ ),
    .Y(\u_ppwm/u_mem/_0014_ ),
    .B1(\u_ppwm/u_mem/_0370_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0876_  (.B1(net514),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0371_ ),
    .VSS(VGND),
    .A1(net424),
    .A2(net298));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0877_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net424),
    .A2(\u_ppwm/u_mem/_0229_ ),
    .Y(\u_ppwm/u_mem/_0015_ ),
    .B1(\u_ppwm/u_mem/_0371_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0878_  (.B1(net514),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0372_ ),
    .VSS(VGND),
    .A1(net434),
    .A2(net561));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0879_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net434),
    .A2(\u_ppwm/u_mem/_0228_ ),
    .Y(\u_ppwm/u_mem/_0016_ ),
    .B1(\u_ppwm/u_mem/_0372_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0880_  (.B1(net516),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0373_ ),
    .VSS(VGND),
    .A1(net433),
    .A2(\u_ppwm/u_mem/memory[10] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0881_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net433),
    .A2(\u_ppwm/u_mem/_0227_ ),
    .Y(\u_ppwm/u_mem/_0017_ ),
    .B1(\u_ppwm/u_mem/_0373_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0882_  (.B1(net515),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0374_ ),
    .VSS(VGND),
    .A1(net433),
    .A2(net280));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0883_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net433),
    .A2(\u_ppwm/u_mem/_0226_ ),
    .Y(\u_ppwm/u_mem/_0018_ ),
    .B1(\u_ppwm/u_mem/_0374_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0884_  (.B1(net515),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0375_ ),
    .VSS(VGND),
    .A1(net432),
    .A2(\u_ppwm/u_mem/memory[12] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0885_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net432),
    .A2(\u_ppwm/u_mem/_0225_ ),
    .Y(\u_ppwm/u_mem/_0019_ ),
    .B1(\u_ppwm/u_mem/_0375_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0886_  (.B1(net513),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0376_ ),
    .VSS(VGND),
    .A1(net432),
    .A2(\u_ppwm/u_mem/memory[13] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0887_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net432),
    .A2(\u_ppwm/u_mem/_0224_ ),
    .Y(\u_ppwm/u_mem/_0020_ ),
    .B1(\u_ppwm/u_mem/_0376_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0888_  (.B1(net513),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0377_ ),
    .VSS(VGND),
    .A1(net423),
    .A2(net275));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0889_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net423),
    .A2(\u_ppwm/u_mem/_0223_ ),
    .Y(\u_ppwm/u_mem/_0021_ ),
    .B1(\u_ppwm/u_mem/_0377_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0890_  (.B1(net514),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0378_ ),
    .VSS(VGND),
    .A1(net434),
    .A2(\u_ppwm/u_mem/memory[15] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0891_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net434),
    .A2(\u_ppwm/u_mem/_0222_ ),
    .Y(\u_ppwm/u_mem/_0022_ ),
    .B1(\u_ppwm/u_mem/_0378_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0892_  (.B1(net516),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0379_ ),
    .VSS(VGND),
    .A1(net435),
    .A2(\u_ppwm/u_mem/memory[16] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0893_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net433),
    .A2(\u_ppwm/u_mem/_0221_ ),
    .Y(\u_ppwm/u_mem/_0023_ ),
    .B1(\u_ppwm/u_mem/_0379_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0894_  (.B1(net515),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0380_ ),
    .VSS(VGND),
    .A1(net436),
    .A2(net543));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0895_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net436),
    .A2(\u_ppwm/u_mem/_0220_ ),
    .Y(\u_ppwm/u_mem/_0024_ ),
    .B1(\u_ppwm/u_mem/_0380_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0896_  (.B1(net515),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0381_ ),
    .VSS(VGND),
    .A1(net436),
    .A2(\u_ppwm/u_mem/memory[18] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0897_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net436),
    .A2(\u_ppwm/u_mem/_0219_ ),
    .Y(\u_ppwm/u_mem/_0025_ ),
    .B1(\u_ppwm/u_mem/_0381_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0898_  (.B1(net511),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0382_ ),
    .VSS(VGND),
    .A1(net432),
    .A2(\u_ppwm/u_mem/memory[19] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0899_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net435),
    .A2(\u_ppwm/u_mem/_0218_ ),
    .Y(\u_ppwm/u_mem/_0026_ ),
    .B1(\u_ppwm/u_mem/_0382_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0900_  (.B1(net513),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0383_ ),
    .VSS(VGND),
    .A1(net432),
    .A2(net331));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0901_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net423),
    .A2(\u_ppwm/u_mem/_0217_ ),
    .Y(\u_ppwm/u_mem/_0027_ ),
    .B1(\u_ppwm/u_mem/_0383_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0902_  (.B1(net513),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0384_ ),
    .VSS(VGND),
    .A1(net424),
    .A2(\u_ppwm/u_mem/memory[21] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0903_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net424),
    .A2(\u_ppwm/u_mem/_0216_ ),
    .Y(\u_ppwm/u_mem/_0028_ ),
    .B1(\u_ppwm/u_mem/_0384_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0904_  (.B1(net514),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0385_ ),
    .VSS(VGND),
    .A1(net424),
    .A2(net282));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0905_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net424),
    .A2(\u_ppwm/u_mem/_0215_ ),
    .Y(\u_ppwm/u_mem/_0029_ ),
    .B1(\u_ppwm/u_mem/_0385_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0906_  (.B1(net513),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0386_ ),
    .VSS(VGND),
    .A1(net434),
    .A2(net524));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0907_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net434),
    .A2(\u_ppwm/u_mem/_0214_ ),
    .Y(\u_ppwm/u_mem/_0030_ ),
    .B1(\u_ppwm/u_mem/_0386_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0908_  (.B1(net515),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0387_ ),
    .VSS(VGND),
    .A1(net436),
    .A2(\u_ppwm/u_mem/memory[24] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0909_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net436),
    .A2(\u_ppwm/u_mem/_0213_ ),
    .Y(\u_ppwm/u_mem/_0031_ ),
    .B1(\u_ppwm/u_mem/_0387_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0910_  (.B1(net515),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0388_ ),
    .VSS(VGND),
    .A1(net436),
    .A2(net262));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0911_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net436),
    .A2(\u_ppwm/u_mem/_0212_ ),
    .Y(\u_ppwm/u_mem/_0032_ ),
    .B1(\u_ppwm/u_mem/_0388_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0912_  (.B1(net511),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0389_ ),
    .VSS(VGND),
    .A1(net435),
    .A2(net336));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0913_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net435),
    .A2(\u_ppwm/u_mem/_0211_ ),
    .Y(\u_ppwm/u_mem/_0033_ ),
    .B1(\u_ppwm/u_mem/_0389_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0914_  (.B1(net512),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0390_ ),
    .VSS(VGND),
    .A1(net426),
    .A2(\u_ppwm/u_mem/memory[27] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0915_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net425),
    .A2(\u_ppwm/u_mem/_0210_ ),
    .Y(\u_ppwm/u_mem/_0034_ ),
    .B1(\u_ppwm/u_mem/_0390_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0916_  (.B1(net512),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0391_ ),
    .VSS(VGND),
    .A1(net425),
    .A2(net288));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0917_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net425),
    .A2(\u_ppwm/u_mem/_0209_ ),
    .Y(\u_ppwm/u_mem/_0035_ ),
    .B1(\u_ppwm/u_mem/_0391_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0918_  (.B1(net512),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0392_ ),
    .VSS(VGND),
    .A1(net426),
    .A2(net329));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0919_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net438),
    .A2(\u_ppwm/u_mem/_0208_ ),
    .Y(\u_ppwm/u_mem/_0036_ ),
    .B1(\u_ppwm/u_mem/_0392_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0920_  (.B1(net510),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0393_ ),
    .VSS(VGND),
    .A1(net426),
    .A2(\u_ppwm/u_mem/memory[30] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0921_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net426),
    .A2(\u_ppwm/u_mem/_0207_ ),
    .Y(\u_ppwm/u_mem/_0037_ ),
    .B1(\u_ppwm/u_mem/_0393_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0922_  (.B1(net510),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0394_ ),
    .VSS(VGND),
    .A1(net427),
    .A2(net324));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0923_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net427),
    .A2(\u_ppwm/u_mem/_0206_ ),
    .Y(\u_ppwm/u_mem/_0038_ ),
    .B1(\u_ppwm/u_mem/_0394_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0924_  (.B1(net502),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0395_ ),
    .VSS(VGND),
    .A1(net419),
    .A2(\u_ppwm/u_mem/memory[32] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0925_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net419),
    .A2(\u_ppwm/u_mem/_0205_ ),
    .Y(\u_ppwm/u_mem/_0039_ ),
    .B1(\u_ppwm/u_mem/_0395_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0926_  (.B1(net502),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0396_ ),
    .VSS(VGND),
    .A1(net417),
    .A2(net226));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0927_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net417),
    .A2(\u_ppwm/u_mem/_0204_ ),
    .Y(\u_ppwm/u_mem/_0040_ ),
    .B1(\u_ppwm/u_mem/_0396_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0928_  (.B1(net504),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0397_ ),
    .VSS(VGND),
    .A1(net417),
    .A2(net314));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0929_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net417),
    .A2(\u_ppwm/u_mem/_0203_ ),
    .Y(\u_ppwm/u_mem/_0041_ ),
    .B1(\u_ppwm/u_mem/_0397_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0930_  (.B1(net512),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0398_ ),
    .VSS(VGND),
    .A1(net425),
    .A2(\u_ppwm/u_mem/memory[35] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0931_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net425),
    .A2(\u_ppwm/u_mem/_0202_ ),
    .Y(\u_ppwm/u_mem/_0042_ ),
    .B1(\u_ppwm/u_mem/_0398_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0932_  (.B1(net512),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0399_ ),
    .VSS(VGND),
    .A1(net425),
    .A2(net220));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0933_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net426),
    .A2(\u_ppwm/u_mem/_0201_ ),
    .Y(\u_ppwm/u_mem/_0043_ ),
    .B1(\u_ppwm/u_mem/_0399_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0934_  (.B1(net510),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0400_ ),
    .VSS(VGND),
    .A1(net426),
    .A2(\u_ppwm/u_mem/memory[37] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0935_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net426),
    .A2(\u_ppwm/u_mem/_0200_ ),
    .Y(\u_ppwm/u_mem/_0044_ ),
    .B1(\u_ppwm/u_mem/_0400_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0936_  (.B1(net502),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0401_ ),
    .VSS(VGND),
    .A1(net426),
    .A2(net320));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0937_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net417),
    .A2(\u_ppwm/u_mem/_0199_ ),
    .Y(\u_ppwm/u_mem/_0045_ ),
    .B1(\u_ppwm/u_mem/_0401_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0938_  (.B1(net502),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0402_ ),
    .VSS(VGND),
    .A1(net421),
    .A2(\u_ppwm/u_mem/memory[39] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0939_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net421),
    .A2(\u_ppwm/u_mem/_0198_ ),
    .Y(\u_ppwm/u_mem/_0046_ ),
    .B1(\u_ppwm/u_mem/_0402_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0940_  (.B1(net502),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0403_ ),
    .VSS(VGND),
    .A1(net417),
    .A2(net273));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0941_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net417),
    .A2(\u_ppwm/u_mem/_0197_ ),
    .Y(\u_ppwm/u_mem/_0047_ ),
    .B1(\u_ppwm/u_mem/_0403_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0942_  (.B1(net510),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0404_ ),
    .VSS(VGND),
    .A1(net427),
    .A2(\u_ppwm/u_mem/memory[41] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0943_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net427),
    .A2(\u_ppwm/u_mem/_0196_ ),
    .Y(\u_ppwm/u_mem/_0048_ ),
    .B1(\u_ppwm/u_mem/_0404_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0944_  (.B1(net511),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0405_ ),
    .VSS(VGND),
    .A1(net429),
    .A2(\u_ppwm/u_mem/memory[42] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0945_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net429),
    .A2(\u_ppwm/u_mem/_0195_ ),
    .Y(\u_ppwm/u_mem/_0049_ ),
    .B1(\u_ppwm/u_mem/_0405_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0946_  (.B1(net511),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0406_ ),
    .VSS(VGND),
    .A1(net429),
    .A2(\u_ppwm/u_mem/memory[43] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0947_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net429),
    .A2(\u_ppwm/u_mem/_0194_ ),
    .Y(\u_ppwm/u_mem/_0050_ ),
    .B1(\u_ppwm/u_mem/_0406_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0948_  (.B1(net511),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0407_ ),
    .VSS(VGND),
    .A1(net430),
    .A2(\u_ppwm/u_mem/memory[44] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0949_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net429),
    .A2(\u_ppwm/u_mem/_0193_ ),
    .Y(\u_ppwm/u_mem/_0051_ ),
    .B1(\u_ppwm/u_mem/_0407_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0950_  (.B1(net510),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0408_ ),
    .VSS(VGND),
    .A1(net427),
    .A2(net278));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0951_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net427),
    .A2(\u_ppwm/u_mem/_0192_ ),
    .Y(\u_ppwm/u_mem/_0052_ ),
    .B1(\u_ppwm/u_mem/_0408_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0952_  (.B1(net510),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0409_ ),
    .VSS(VGND),
    .A1(net427),
    .A2(\u_ppwm/u_mem/memory[46] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0953_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net428),
    .A2(\u_ppwm/u_mem/_0191_ ),
    .Y(\u_ppwm/u_mem/_0053_ ),
    .B1(\u_ppwm/u_mem/_0409_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0954_  (.B1(net502),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0410_ ),
    .VSS(VGND),
    .A1(net419),
    .A2(\u_ppwm/u_mem/memory[47] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0955_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net419),
    .A2(\u_ppwm/u_mem/_0190_ ),
    .Y(\u_ppwm/u_mem/_0054_ ),
    .B1(\u_ppwm/u_mem/_0410_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0956_  (.B1(net502),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0411_ ),
    .VSS(VGND),
    .A1(net419),
    .A2(net240));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0957_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net419),
    .A2(\u_ppwm/u_mem/_0189_ ),
    .Y(\u_ppwm/u_mem/_0055_ ),
    .B1(\u_ppwm/u_mem/_0411_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0958_  (.B1(net510),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0412_ ),
    .VSS(VGND),
    .A1(net429),
    .A2(net309));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0959_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net429),
    .A2(\u_ppwm/u_mem/_0188_ ),
    .Y(\u_ppwm/u_mem/_0056_ ),
    .B1(\u_ppwm/u_mem/_0412_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0960_  (.B1(net511),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0413_ ),
    .VSS(VGND),
    .A1(net430),
    .A2(\u_ppwm/u_mem/memory[50] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0961_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net430),
    .A2(\u_ppwm/u_mem/_0187_ ),
    .Y(\u_ppwm/u_mem/_0057_ ),
    .B1(\u_ppwm/u_mem/_0413_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0962_  (.B1(net512),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0414_ ),
    .VSS(VGND),
    .A1(net429),
    .A2(net245));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0963_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net430),
    .A2(\u_ppwm/u_mem/_0186_ ),
    .Y(\u_ppwm/u_mem/_0058_ ),
    .B1(\u_ppwm/u_mem/_0414_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0964_  (.B1(net510),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0415_ ),
    .VSS(VGND),
    .A1(net427),
    .A2(net536));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0965_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net428),
    .A2(\u_ppwm/u_mem/_0185_ ),
    .Y(\u_ppwm/u_mem/_0059_ ),
    .B1(\u_ppwm/u_mem/_0415_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0966_  (.B1(net511),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0416_ ),
    .VSS(VGND),
    .A1(net428),
    .A2(\u_ppwm/u_mem/memory[53] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0967_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net428),
    .A2(\u_ppwm/u_mem/_0184_ ),
    .Y(\u_ppwm/u_mem/_0060_ ),
    .B1(\u_ppwm/u_mem/_0416_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0968_  (.B1(net502),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0417_ ),
    .VSS(VGND),
    .A1(net420),
    .A2(net271));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0969_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net420),
    .A2(\u_ppwm/u_mem/_0183_ ),
    .Y(\u_ppwm/u_mem/_0061_ ),
    .B1(\u_ppwm/u_mem/_0417_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0970_  (.B1(net503),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0418_ ),
    .VSS(VGND),
    .A1(net419),
    .A2(\u_ppwm/u_mem/memory[55] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0971_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net419),
    .A2(\u_ppwm/u_mem/_0182_ ),
    .Y(\u_ppwm/u_mem/_0062_ ),
    .B1(\u_ppwm/u_mem/_0418_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0972_  (.B1(net503),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0419_ ),
    .VSS(VGND),
    .A1(net420),
    .A2(net286));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0973_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net420),
    .A2(\u_ppwm/u_mem/_0181_ ),
    .Y(\u_ppwm/u_mem/_0063_ ),
    .B1(\u_ppwm/u_mem/_0419_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0974_  (.B1(net498),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0420_ ),
    .VSS(VGND),
    .A1(net415),
    .A2(\u_ppwm/u_mem/memory[57] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0975_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net415),
    .A2(\u_ppwm/u_mem/_0180_ ),
    .Y(\u_ppwm/u_mem/_0064_ ),
    .B1(\u_ppwm/u_mem/_0420_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0976_  (.B1(net496),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0421_ ),
    .VSS(VGND),
    .A1(net412),
    .A2(\u_ppwm/u_mem/memory[58] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0977_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net413),
    .A2(\u_ppwm/u_mem/_0179_ ),
    .Y(\u_ppwm/u_mem/_0065_ ),
    .B1(\u_ppwm/u_mem/_0421_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0978_  (.B1(net497),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0422_ ),
    .VSS(VGND),
    .A1(net413),
    .A2(net224));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0979_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net413),
    .A2(\u_ppwm/u_mem/_0178_ ),
    .Y(\u_ppwm/u_mem/_0066_ ),
    .B1(\u_ppwm/u_mem/_0422_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0980_  (.B1(net496),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0423_ ),
    .VSS(VGND),
    .A1(net412),
    .A2(net264));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0981_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net409),
    .A2(\u_ppwm/u_mem/_0177_ ),
    .Y(\u_ppwm/u_mem/_0067_ ),
    .B1(\u_ppwm/u_mem/_0423_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0982_  (.B1(net496),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0424_ ),
    .VSS(VGND),
    .A1(net409),
    .A2(net306));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0983_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net409),
    .A2(\u_ppwm/u_mem/_0176_ ),
    .Y(\u_ppwm/u_mem/_0068_ ),
    .B1(\u_ppwm/u_mem/_0424_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0984_  (.B1(net498),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0425_ ),
    .VSS(VGND),
    .A1(net415),
    .A2(\u_ppwm/u_mem/memory[62] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0985_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net415),
    .A2(\u_ppwm/u_mem/_0175_ ),
    .Y(\u_ppwm/u_mem/_0069_ ),
    .B1(\u_ppwm/u_mem/_0425_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0986_  (.B1(net503),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0426_ ),
    .VSS(VGND),
    .A1(net420),
    .A2(\u_ppwm/u_mem/memory[63] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0987_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net420),
    .A2(\u_ppwm/u_mem/_0174_ ),
    .Y(\u_ppwm/u_mem/_0070_ ),
    .B1(\u_ppwm/u_mem/_0426_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0988_  (.B1(net498),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0427_ ),
    .VSS(VGND),
    .A1(net415),
    .A2(net251));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0989_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net416),
    .A2(\u_ppwm/u_mem/_0173_ ),
    .Y(\u_ppwm/u_mem/_0071_ ),
    .B1(\u_ppwm/u_mem/_0427_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0990_  (.B1(net497),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0428_ ),
    .VSS(VGND),
    .A1(net413),
    .A2(\u_ppwm/u_mem/memory[65] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0991_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net413),
    .A2(\u_ppwm/u_mem/_0172_ ),
    .Y(\u_ppwm/u_mem/_0072_ ),
    .B1(\u_ppwm/u_mem/_0428_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0992_  (.B1(net497),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0429_ ),
    .VSS(VGND),
    .A1(net413),
    .A2(net228));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0993_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net413),
    .A2(\u_ppwm/u_mem/_0171_ ),
    .Y(\u_ppwm/u_mem/_0073_ ),
    .B1(\u_ppwm/u_mem/_0429_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0994_  (.B1(net496),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0430_ ),
    .VSS(VGND),
    .A1(net412),
    .A2(net292));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0995_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net409),
    .A2(\u_ppwm/u_mem/_0170_ ),
    .Y(\u_ppwm/u_mem/_0074_ ),
    .B1(\u_ppwm/u_mem/_0430_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0996_  (.B1(net496),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0431_ ),
    .VSS(VGND),
    .A1(net410),
    .A2(net297));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0997_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net410),
    .A2(\u_ppwm/u_mem/_0169_ ),
    .Y(\u_ppwm/u_mem/_0075_ ),
    .B1(\u_ppwm/u_mem/_0431_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0998_  (.B1(net498),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0432_ ),
    .VSS(VGND),
    .A1(net411),
    .A2(\u_ppwm/u_mem/memory[69] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0999_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net411),
    .A2(\u_ppwm/u_mem/_0168_ ),
    .Y(\u_ppwm/u_mem/_0076_ ),
    .B1(\u_ppwm/u_mem/_0432_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1000_  (.B1(net498),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0433_ ),
    .VSS(VGND),
    .A1(net414),
    .A2(\u_ppwm/u_mem/memory[70] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1001_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net414),
    .A2(\u_ppwm/u_mem/_0167_ ),
    .Y(\u_ppwm/u_mem/_0077_ ),
    .B1(\u_ppwm/u_mem/_0433_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1002_  (.B1(net498),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0434_ ),
    .VSS(VGND),
    .A1(net415),
    .A2(\u_ppwm/u_mem/memory[71] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1003_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net415),
    .A2(\u_ppwm/u_mem/_0166_ ),
    .Y(\u_ppwm/u_mem/_0078_ ),
    .B1(\u_ppwm/u_mem/_0434_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1004_  (.B1(net499),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0435_ ),
    .VSS(VGND),
    .A1(net414),
    .A2(\u_ppwm/u_mem/memory[72] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1005_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net412),
    .A2(\u_ppwm/u_mem/_0165_ ),
    .Y(\u_ppwm/u_mem/_0079_ ),
    .B1(\u_ppwm/u_mem/_0435_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1006_  (.B1(net497),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0436_ ),
    .VSS(VGND),
    .A1(net412),
    .A2(net234));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1007_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net412),
    .A2(\u_ppwm/u_mem/_0164_ ),
    .Y(\u_ppwm/u_mem/_0080_ ),
    .B1(\u_ppwm/u_mem/_0436_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1008_  (.B1(net496),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0437_ ),
    .VSS(VGND),
    .A1(net409),
    .A2(net244));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1009_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net409),
    .A2(\u_ppwm/u_mem/_0163_ ),
    .Y(\u_ppwm/u_mem/_0081_ ),
    .B1(\u_ppwm/u_mem/_0437_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1010_  (.B1(net495),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0438_ ),
    .VSS(VGND),
    .A1(net410),
    .A2(\u_ppwm/u_mem/memory[75] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1011_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net410),
    .A2(\u_ppwm/u_mem/_0162_ ),
    .Y(\u_ppwm/u_mem/_0082_ ),
    .B1(\u_ppwm/u_mem/_0438_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1012_  (.B1(net494),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0439_ ),
    .VSS(VGND),
    .A1(net411),
    .A2(net345));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1013_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net411),
    .A2(\u_ppwm/u_mem/_0161_ ),
    .Y(\u_ppwm/u_mem/_0083_ ),
    .B1(\u_ppwm/u_mem/_0439_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1014_  (.B1(net498),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0440_ ),
    .VSS(VGND),
    .A1(net411),
    .A2(\u_ppwm/u_mem/memory[77] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1015_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net414),
    .A2(\u_ppwm/u_mem/_0160_ ),
    .Y(\u_ppwm/u_mem/_0084_ ),
    .B1(\u_ppwm/u_mem/_0440_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1016_  (.B1(net498),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0441_ ),
    .VSS(VGND),
    .A1(net414),
    .A2(\u_ppwm/u_mem/memory[78] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1017_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net414),
    .A2(\u_ppwm/u_mem/_0159_ ),
    .Y(\u_ppwm/u_mem/_0085_ ),
    .B1(\u_ppwm/u_mem/_0441_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1018_  (.B1(net499),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0442_ ),
    .VSS(VGND),
    .A1(net414),
    .A2(\u_ppwm/u_mem/memory[79] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1019_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net414),
    .A2(\u_ppwm/u_mem/_0158_ ),
    .Y(\u_ppwm/u_mem/_0086_ ),
    .B1(\u_ppwm/u_mem/_0442_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1020_  (.B1(net496),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0443_ ),
    .VSS(VGND),
    .A1(net412),
    .A2(net236));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1021_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net412),
    .A2(\u_ppwm/u_mem/_0157_ ),
    .Y(\u_ppwm/u_mem/_0087_ ),
    .B1(\u_ppwm/u_mem/_0443_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1022_  (.B1(net496),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0444_ ),
    .VSS(VGND),
    .A1(net409),
    .A2(net319));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1023_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net409),
    .A2(\u_ppwm/u_mem/_0156_ ),
    .Y(\u_ppwm/u_mem/_0088_ ),
    .B1(\u_ppwm/u_mem/_0444_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1024_  (.B1(net495),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0445_ ),
    .VSS(VGND),
    .A1(net410),
    .A2(\u_ppwm/u_mem/memory[82] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1025_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net410),
    .A2(\u_ppwm/u_mem/_0155_ ),
    .Y(\u_ppwm/u_mem/_0089_ ),
    .B1(\u_ppwm/u_mem/_0445_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1026_  (.B1(net494),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0446_ ),
    .VSS(VGND),
    .A1(net404),
    .A2(net326));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1027_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net404),
    .A2(\u_ppwm/u_mem/_0154_ ),
    .Y(\u_ppwm/u_mem/_0090_ ),
    .B1(\u_ppwm/u_mem/_0446_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1028_  (.B1(net495),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0447_ ),
    .VSS(VGND),
    .A1(net405),
    .A2(\u_ppwm/u_mem/memory[84] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1029_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net405),
    .A2(\u_ppwm/u_mem/_0153_ ),
    .Y(\u_ppwm/u_mem/_0091_ ),
    .B1(\u_ppwm/u_mem/_0447_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1030_  (.B1(net495),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0448_ ),
    .VSS(VGND),
    .A1(net411),
    .A2(net538));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1031_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net411),
    .A2(\u_ppwm/u_mem/_0152_ ),
    .Y(\u_ppwm/u_mem/_0092_ ),
    .B1(\u_ppwm/u_mem/_0448_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1032_  (.B1(net503),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0449_ ),
    .VSS(VGND),
    .A1(net418),
    .A2(\u_ppwm/u_mem/memory[86] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1033_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net418),
    .A2(\u_ppwm/u_mem/_0151_ ),
    .Y(\u_ppwm/u_mem/_0093_ ),
    .B1(\u_ppwm/u_mem/_0449_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1034_  (.B1(net501),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0450_ ),
    .VSS(VGND),
    .A1(net418),
    .A2(net230));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1035_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net418),
    .A2(\u_ppwm/u_mem/_0150_ ),
    .Y(\u_ppwm/u_mem/_0094_ ),
    .B1(\u_ppwm/u_mem/_0450_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1036_  (.B1(net501),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0451_ ),
    .VSS(VGND),
    .A1(net407),
    .A2(\u_ppwm/u_mem/memory[88] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1037_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net407),
    .A2(\u_ppwm/u_mem/_0149_ ),
    .Y(\u_ppwm/u_mem/_0095_ ),
    .B1(\u_ppwm/u_mem/_0451_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1038_  (.B1(net501),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0452_ ),
    .VSS(VGND),
    .A1(net407),
    .A2(net232));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1039_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net407),
    .A2(\u_ppwm/u_mem/_0148_ ),
    .Y(\u_ppwm/u_mem/_0096_ ),
    .B1(\u_ppwm/u_mem/_0452_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1040_  (.B1(net500),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0453_ ),
    .VSS(VGND),
    .A1(net405),
    .A2(\u_ppwm/u_mem/memory[90] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1041_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net405),
    .A2(\u_ppwm/u_mem/_0147_ ),
    .Y(\u_ppwm/u_mem/_0097_ ),
    .B1(\u_ppwm/u_mem/_0453_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1042_  (.B1(net495),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0454_ ),
    .VSS(VGND),
    .A1(net405),
    .A2(net205));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1043_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net405),
    .A2(\u_ppwm/u_mem/_0146_ ),
    .Y(\u_ppwm/u_mem/_0098_ ),
    .B1(\u_ppwm/u_mem/_0454_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1044_  (.B1(net495),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0455_ ),
    .VSS(VGND),
    .A1(net405),
    .A2(net526));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1045_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net407),
    .A2(\u_ppwm/u_mem/_0145_ ),
    .Y(\u_ppwm/u_mem/_0099_ ),
    .B1(\u_ppwm/u_mem/_0455_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1046_  (.B1(net503),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0456_ ),
    .VSS(VGND),
    .A1(net418),
    .A2(\u_ppwm/u_mem/memory[93] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1047_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net418),
    .A2(\u_ppwm/u_mem/_0144_ ),
    .Y(\u_ppwm/u_mem/_0100_ ),
    .B1(\u_ppwm/u_mem/_0456_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1048_  (.B1(net501),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0457_ ),
    .VSS(VGND),
    .A1(net418),
    .A2(\u_ppwm/u_mem/memory[94] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1049_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net417),
    .A2(\u_ppwm/u_mem/_0143_ ),
    .Y(\u_ppwm/u_mem/_0101_ ),
    .B1(\u_ppwm/u_mem/_0457_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1050_  (.B1(net501),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0458_ ),
    .VSS(VGND),
    .A1(net408),
    .A2(\u_ppwm/u_mem/memory[95] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1051_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net407),
    .A2(\u_ppwm/u_mem/_0142_ ),
    .Y(\u_ppwm/u_mem/_0102_ ),
    .B1(\u_ppwm/u_mem/_0458_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1052_  (.B1(net501),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0459_ ),
    .VSS(VGND),
    .A1(net407),
    .A2(net213));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1053_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net407),
    .A2(\u_ppwm/u_mem/_0141_ ),
    .Y(\u_ppwm/u_mem/_0103_ ),
    .B1(\u_ppwm/u_mem/_0459_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1054_  (.B1(net501),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0460_ ),
    .VSS(VGND),
    .A1(net408),
    .A2(\u_ppwm/u_mem/memory[97] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1055_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net408),
    .A2(\u_ppwm/u_mem/_0140_ ),
    .Y(\u_ppwm/u_mem/_0104_ ),
    .B1(\u_ppwm/u_mem/_0460_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1056_  (.B1(net488),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0461_ ),
    .VSS(VGND),
    .A1(net402),
    .A2(\u_ppwm/u_mem/memory[98] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1057_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net402),
    .A2(\u_ppwm/u_mem/_0139_ ),
    .Y(\u_ppwm/u_mem/_0105_ ),
    .B1(\u_ppwm/u_mem/_0461_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1058_  (.B1(net488),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0462_ ),
    .VSS(VGND),
    .A1(net402),
    .A2(\u_ppwm/u_mem/memory[99] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1059_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net402),
    .A2(\u_ppwm/u_mem/_0138_ ),
    .Y(\u_ppwm/u_mem/_0106_ ),
    .B1(\u_ppwm/u_mem/_0462_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1060_  (.B1(net500),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0463_ ),
    .VSS(VGND),
    .A1(net406),
    .A2(\u_ppwm/u_mem/memory[100] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1061_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net403),
    .A2(\u_ppwm/u_mem/_0137_ ),
    .Y(\u_ppwm/u_mem/_0107_ ),
    .B1(\u_ppwm/u_mem/_0463_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1062_  (.B1(net494),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0464_ ),
    .VSS(VGND),
    .A1(net403),
    .A2(net253));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1063_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net403),
    .A2(\u_ppwm/u_mem/_0136_ ),
    .Y(\u_ppwm/u_mem/_0108_ ),
    .B1(\u_ppwm/u_mem/_0464_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1064_  (.B1(net494),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0465_ ),
    .VSS(VGND),
    .A1(net403),
    .A2(net318));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1065_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net403),
    .A2(\u_ppwm/u_mem/_0135_ ),
    .Y(\u_ppwm/u_mem/_0109_ ),
    .B1(\u_ppwm/u_mem/_0465_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1066_  (.B1(net494),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0466_ ),
    .VSS(VGND),
    .A1(net401),
    .A2(net528));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1067_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net401),
    .A2(\u_ppwm/u_mem/_0134_ ),
    .Y(\u_ppwm/u_mem/_0110_ ),
    .B1(\u_ppwm/u_mem/_0466_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1068_  (.B1(net488),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0467_ ),
    .VSS(VGND),
    .A1(net401),
    .A2(\u_ppwm/u_mem/memory[104] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1069_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net401),
    .A2(\u_ppwm/u_mem/_0133_ ),
    .Y(\u_ppwm/u_mem/_0111_ ),
    .B1(\u_ppwm/u_mem/_0467_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1070_  (.B1(net493),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0468_ ),
    .VSS(VGND),
    .A1(net406),
    .A2(\u_ppwm/u_mem/memory[105] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1071_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net402),
    .A2(\u_ppwm/u_mem/_0132_ ),
    .Y(\u_ppwm/u_mem/_0112_ ),
    .B1(\u_ppwm/u_mem/_0468_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1072_  (.B1(net500),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0469_ ),
    .VSS(VGND),
    .A1(net402),
    .A2(\u_ppwm/u_mem/memory[106] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1073_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net406),
    .A2(\u_ppwm/u_mem/_0131_ ),
    .Y(\u_ppwm/u_mem/_0113_ ),
    .B1(\u_ppwm/u_mem/_0469_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1074_  (.B1(net494),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0470_ ),
    .VSS(VGND),
    .A1(net403),
    .A2(\u_ppwm/u_mem/memory[107] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1075_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net404),
    .A2(\u_ppwm/u_mem/_0130_ ),
    .Y(\u_ppwm/u_mem/_0114_ ),
    .B1(\u_ppwm/u_mem/_0470_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1076_  (.B1(net495),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0471_ ),
    .VSS(VGND),
    .A1(net404),
    .A2(net222));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1077_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net404),
    .A2(\u_ppwm/u_mem/_0129_ ),
    .Y(\u_ppwm/u_mem/_0115_ ),
    .B1(\u_ppwm/u_mem/_0471_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1078_  (.B1(net494),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0472_ ),
    .VSS(VGND),
    .A1(net403),
    .A2(\u_ppwm/u_mem/_0001_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1079_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net403),
    .A2(\u_ppwm/u_mem/_0128_ ),
    .Y(\u_ppwm/u_mem/_0116_ ),
    .B1(\u_ppwm/u_mem/_0472_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1080_  (.B1(net494),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0473_ ),
    .VSS(VGND),
    .A1(net400),
    .A2(net295));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1081_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0126_ ),
    .A2(net400),
    .Y(\u_ppwm/u_mem/_0117_ ),
    .B1(\u_ppwm/u_mem/_0473_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1082_  (.B1(net488),
    .VDD(VPWR),
    .Y(\u_ppwm/u_mem/_0474_ ),
    .VSS(VGND),
    .A1(net535),
    .A2(net401));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1083_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_mem/_0127_ ),
    .A2(net400),
    .Y(\u_ppwm/u_mem/_0118_ ),
    .B1(\u_ppwm/u_mem/_0474_ ));
 sg13g2_nand2b_2 \u_ppwm/u_mem/_1084_  (.Y(\u_ppwm/u_mem/_0475_ ),
    .B(net333),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net400));
 sg13g2_nand2_2 \u_ppwm/u_mem/_1085_  (.Y(\u_ppwm/u_mem/_0476_ ),
    .A(net488),
    .B(\u_ppwm/u_mem/_0475_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1086_  (.A(net617),
    .B(net400),
    .Y(\u_ppwm/u_mem/_0477_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_mem/_1087_  (.A(net617),
    .B(net400),
    .X(\u_ppwm/u_mem/_0478_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1088_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(\u_ppwm/u_mem/_0477_ ),
    .C(\u_ppwm/u_mem/_0478_ ),
    .Y(\u_ppwm/u_mem/_0119_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1089_  (.A(net638),
    .B(\u_ppwm/u_mem/_0478_ ),
    .Y(\u_ppwm/u_mem/_0479_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_mem/_1090_  (.A(net638),
    .B(\u_ppwm/u_mem/_0478_ ),
    .X(\u_ppwm/u_mem/_0480_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1091_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(\u_ppwm/u_mem/_0479_ ),
    .C(\u_ppwm/u_mem/_0480_ ),
    .Y(\u_ppwm/u_mem/_0120_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1092_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net611),
    .A2(\u_ppwm/u_mem/_0475_ ),
    .Y(\u_ppwm/u_mem/_0481_ ),
    .B1(\u_ppwm/u_mem/_0480_ ));
 sg13g2_and4_1 \u_ppwm/u_mem/_1093_  (.A(net611),
    .B(net691),
    .C(net624),
    .D(net400),
    .X(\u_ppwm/u_mem/_0482_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1094_  (.A(\u_ppwm/u_mem/_0238_ ),
    .B(net612),
    .C(\u_ppwm/u_mem/_0482_ ),
    .Y(\u_ppwm/u_mem/_0121_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1095_  (.A(net606),
    .B(\u_ppwm/u_mem/_0482_ ),
    .Y(\u_ppwm/u_mem/_0483_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_mem/_1096_  (.A(net606),
    .B(\u_ppwm/u_mem/_0482_ ),
    .X(\u_ppwm/u_mem/_0484_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1097_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(net607),
    .C(\u_ppwm/u_mem/_0484_ ),
    .Y(\u_ppwm/u_mem/_0122_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1098_  (.A(net618),
    .B(\u_ppwm/u_mem/_0484_ ),
    .Y(\u_ppwm/u_mem/_0485_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 \u_ppwm/u_mem/_1099_  (.X(\u_ppwm/u_mem/_0486_ ),
    .A(net618),
    .B(net606),
    .C(\u_ppwm/u_mem/_0482_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1100_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(\u_ppwm/u_mem/_0485_ ),
    .C(\u_ppwm/u_mem/_0486_ ),
    .Y(\u_ppwm/u_mem/_0123_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1101_  (.A(net587),
    .B(\u_ppwm/u_mem/_0486_ ),
    .Y(\u_ppwm/u_mem/_0487_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 \u_ppwm/u_mem/_1102_  (.A(net587),
    .B(\u_ppwm/u_mem/bit_count[4] ),
    .C(\u_ppwm/u_mem/bit_count[3] ),
    .D(\u_ppwm/u_mem/_0482_ ),
    .X(\u_ppwm/u_mem/_0488_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1103_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(net588),
    .C(\u_ppwm/u_mem/_0488_ ),
    .Y(\u_ppwm/u_mem/_0124_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1104_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net565),
    .A2(\u_ppwm/u_mem/_0475_ ),
    .Y(\u_ppwm/u_mem/_0489_ ),
    .B1(\u_ppwm/u_mem/_0488_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1105_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net565),
    .A2(\u_ppwm/u_mem/_0488_ ),
    .Y(\u_ppwm/u_mem/_0490_ ),
    .B1(\u_ppwm/u_mem/_0238_ ));
 sg13g2_nor2b_1 \u_ppwm/u_mem/_1106_  (.A(net566),
    .B_N(\u_ppwm/u_mem/_0490_ ),
    .Y(\u_ppwm/u_mem/_0125_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1107_  (.RESET_B(net174),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net598),
    .Q(\u_ppwm/u_mem/memory[0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1108_  (.RESET_B(net146),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net578),
    .Q(\u_ppwm/u_mem/memory[1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1109_  (.RESET_B(net144),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net342),
    .Q(\u_ppwm/u_mem/memory[2] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1110_  (.RESET_B(net142),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net243),
    .Q(\u_ppwm/u_mem/memory[3] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1111_  (.RESET_B(net140),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0011_ ),
    .Q(\u_ppwm/u_mem/memory[4] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1112_  (.RESET_B(net138),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0012_ ),
    .Q(\u_ppwm/u_mem/memory[5] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1113_  (.RESET_B(net136),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net285),
    .Q(\u_ppwm/u_mem/memory[6] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1114_  (.RESET_B(net134),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0014_ ),
    .Q(\u_ppwm/u_mem/memory[7] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1115_  (.RESET_B(net132),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net562),
    .Q(\u_ppwm/u_mem/memory[8] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1116_  (.RESET_B(net130),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0016_ ),
    .Q(\u_ppwm/u_mem/memory[9] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1117_  (.RESET_B(net128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net281),
    .Q(\u_ppwm/u_mem/memory[10] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1118_  (.RESET_B(net126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0018_ ),
    .Q(\u_ppwm/u_mem/memory[11] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1119_  (.RESET_B(net124),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net294),
    .Q(\u_ppwm/u_mem/memory[12] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1120_  (.RESET_B(net122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net276),
    .Q(\u_ppwm/u_mem/memory[13] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1121_  (.RESET_B(net120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0021_ ),
    .Q(\u_ppwm/u_mem/memory[14] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1122_  (.RESET_B(net118),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net552),
    .Q(\u_ppwm/u_mem/memory[15] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1123_  (.RESET_B(net116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net544),
    .Q(\u_ppwm/u_mem/memory[16] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1124_  (.RESET_B(net114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0024_ ),
    .Q(\u_ppwm/u_mem/memory[17] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1125_  (.RESET_B(net112),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net530),
    .Q(\u_ppwm/u_mem/memory[18] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1126_  (.RESET_B(net110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net332),
    .Q(\u_ppwm/u_mem/memory[19] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1127_  (.RESET_B(net108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0027_ ),
    .Q(\u_ppwm/u_mem/memory[20] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1128_  (.RESET_B(net106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net283),
    .Q(\u_ppwm/u_mem/memory[21] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1129_  (.RESET_B(net104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net525),
    .Q(\u_ppwm/u_mem/memory[22] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1130_  (.RESET_B(net102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0030_ ),
    .Q(\u_ppwm/u_mem/memory[23] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1131_  (.RESET_B(net100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net263),
    .Q(\u_ppwm/u_mem/memory[24] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1132_  (.RESET_B(net98),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0032_ ),
    .Q(\u_ppwm/u_mem/memory[25] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1133_  (.RESET_B(net96),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0033_ ),
    .Q(\u_ppwm/u_mem/memory[26] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1134_  (.RESET_B(net94),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net289),
    .Q(\u_ppwm/u_mem/memory[27] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1135_  (.RESET_B(net92),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net330),
    .Q(\u_ppwm/u_mem/memory[28] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1136_  (.RESET_B(net90),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net555),
    .Q(\u_ppwm/u_mem/memory[29] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1137_  (.RESET_B(net88),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net325),
    .Q(\u_ppwm/u_mem/memory[30] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1138_  (.RESET_B(net86),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0038_ ),
    .Q(\u_ppwm/u_mem/memory[31] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1139_  (.RESET_B(net84),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net227),
    .Q(\u_ppwm/u_mem/memory[32] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1140_  (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0040_ ),
    .Q(\u_ppwm/u_mem/memory[33] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1141_  (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0041_ ),
    .Q(\u_ppwm/u_mem/memory[34] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1142_  (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net221),
    .Q(\u_ppwm/u_mem/memory[35] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1143_  (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net338),
    .Q(\u_ppwm/u_mem/memory[36] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1144_  (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net321),
    .Q(\u_ppwm/u_mem/memory[37] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1145_  (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0045_ ),
    .Q(\u_ppwm/u_mem/memory[38] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1146_  (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net274),
    .Q(\u_ppwm/u_mem/memory[39] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1147_  (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0047_ ),
    .Q(\u_ppwm/u_mem/memory[40] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1148_  (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net557),
    .Q(\u_ppwm/u_mem/memory[41] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1149_  (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net523),
    .Q(\u_ppwm/u_mem/memory[42] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1150_  (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net311),
    .Q(\u_ppwm/u_mem/memory[43] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1151_  (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net279),
    .Q(\u_ppwm/u_mem/memory[44] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1152_  (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0052_ ),
    .Q(\u_ppwm/u_mem/memory[45] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1153_  (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net270),
    .Q(\u_ppwm/u_mem/memory[46] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1154_  (.RESET_B(net173),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net241),
    .Q(\u_ppwm/u_mem/memory[47] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1155_  (.RESET_B(net171),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0055_ ),
    .Q(\u_ppwm/u_mem/memory[48] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1156_  (.RESET_B(net169),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0056_ ),
    .Q(\u_ppwm/u_mem/memory[49] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1157_  (.RESET_B(net167),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net246),
    .Q(\u_ppwm/u_mem/memory[50] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1158_  (.RESET_B(net165),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0058_ ),
    .Q(\u_ppwm/u_mem/memory[51] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1159_  (.RESET_B(net163),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0059_ ),
    .Q(\u_ppwm/u_mem/memory[52] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1160_  (.RESET_B(net161),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net272),
    .Q(\u_ppwm/u_mem/memory[53] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1161_  (.RESET_B(net159),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0061_ ),
    .Q(\u_ppwm/u_mem/memory[54] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1162_  (.RESET_B(net157),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net287),
    .Q(\u_ppwm/u_mem/memory[55] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1163_  (.RESET_B(net155),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0063_ ),
    .Q(\u_ppwm/u_mem/memory[56] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1164_  (.RESET_B(net153),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net316),
    .Q(\u_ppwm/u_mem/memory[57] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1165_  (.RESET_B(net151),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net225),
    .Q(\u_ppwm/u_mem/memory[58] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1166_  (.RESET_B(net149),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0066_ ),
    .Q(\u_ppwm/u_mem/memory[59] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1167_  (.RESET_B(net147),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0067_ ),
    .Q(\u_ppwm/u_mem/memory[60] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1168_  (.RESET_B(net143),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0068_ ),
    .Q(\u_ppwm/u_mem/memory[61] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1169_  (.RESET_B(net139),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net268),
    .Q(\u_ppwm/u_mem/memory[62] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1170_  (.RESET_B(net135),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net252),
    .Q(\u_ppwm/u_mem/memory[63] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1171_  (.RESET_B(net131),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net304),
    .Q(\u_ppwm/u_mem/memory[64] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1172_  (.RESET_B(net127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net229),
    .Q(\u_ppwm/u_mem/memory[65] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1173_  (.RESET_B(net123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0073_ ),
    .Q(\u_ppwm/u_mem/memory[66] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1174_  (.RESET_B(net119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0074_ ),
    .Q(\u_ppwm/u_mem/memory[67] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1175_  (.RESET_B(net115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0075_ ),
    .Q(\u_ppwm/u_mem/memory[68] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1176_  (.RESET_B(net111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net519),
    .Q(\u_ppwm/u_mem/memory[69] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1177_  (.RESET_B(net107),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net266),
    .Q(\u_ppwm/u_mem/memory[70] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1178_  (.RESET_B(net103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net256),
    .Q(\u_ppwm/u_mem/memory[71] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1179_  (.RESET_B(net99),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net235),
    .Q(\u_ppwm/u_mem/memory[72] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1180_  (.RESET_B(net95),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0080_ ),
    .Q(\u_ppwm/u_mem/memory[73] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1181_  (.RESET_B(net91),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0081_ ),
    .Q(\u_ppwm/u_mem/memory[74] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1182_  (.RESET_B(net87),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net346),
    .Q(\u_ppwm/u_mem/memory[75] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1183_  (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net584),
    .Q(\u_ppwm/u_mem/memory[76] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1184_  (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net323),
    .Q(\u_ppwm/u_mem/memory[77] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1185_  (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net250),
    .Q(\u_ppwm/u_mem/memory[78] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1186_  (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net237),
    .Q(\u_ppwm/u_mem/memory[79] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1187_  (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0087_ ),
    .Q(\u_ppwm/u_mem/memory[80] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1188_  (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0088_ ),
    .Q(\u_ppwm/u_mem/memory[81] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1189_  (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net327),
    .Q(\u_ppwm/u_mem/memory[82] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1190_  (.RESET_B(net55),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0090_ ),
    .Q(\u_ppwm/u_mem/memory[83] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1191_  (.RESET_B(net170),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net539),
    .Q(\u_ppwm/u_mem/memory[84] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1192_  (.RESET_B(net166),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net569),
    .Q(\u_ppwm/u_mem/memory[85] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1193_  (.RESET_B(net162),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net231),
    .Q(\u_ppwm/u_mem/memory[86] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1194_  (.RESET_B(net158),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0094_ ),
    .Q(\u_ppwm/u_mem/memory[87] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1195_  (.RESET_B(net154),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net233),
    .Q(\u_ppwm/u_mem/memory[88] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1196_  (.RESET_B(net150),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0096_ ),
    .Q(\u_ppwm/u_mem/memory[89] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1197_  (.RESET_B(net145),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net206),
    .Q(\u_ppwm/u_mem/memory[90] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1198_  (.RESET_B(net137),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0098_ ),
    .Q(\u_ppwm/u_mem/memory[91] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1199_  (.RESET_B(net129),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0099_ ),
    .Q(\u_ppwm/u_mem/memory[92] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1200_  (.RESET_B(net121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net521),
    .Q(\u_ppwm/u_mem/memory[93] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1201_  (.RESET_B(net113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net340),
    .Q(\u_ppwm/u_mem/memory[94] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1202_  (.RESET_B(net105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net214),
    .Q(\u_ppwm/u_mem/memory[95] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1203_  (.RESET_B(net97),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0103_ ),
    .Q(\u_ppwm/u_mem/memory[96] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1204_  (.RESET_B(net89),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net313),
    .Q(\u_ppwm/u_mem/memory[97] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1205_  (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net302),
    .Q(\u_ppwm/u_mem/memory[98] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1206_  (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net259),
    .Q(\u_ppwm/u_mem/memory[99] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1207_  (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net254),
    .Q(\u_ppwm/u_mem/memory[100] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1208_  (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0108_ ),
    .Q(\u_ppwm/u_mem/memory[101] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1209_  (.RESET_B(net168),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0109_ ),
    .Q(\u_ppwm/u_mem/memory[102] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1210_  (.RESET_B(net160),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0110_ ),
    .Q(\u_ppwm/u_mem/memory[103] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1211_  (.RESET_B(net152),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net344),
    .Q(\u_ppwm/u_mem/memory[104] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1212_  (.RESET_B(net141),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net308),
    .Q(\u_ppwm/u_mem/memory[105] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1213_  (.RESET_B(net125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net291),
    .Q(\u_ppwm/u_mem/memory[106] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1214_  (.RESET_B(net109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net223),
    .Q(\u_ppwm/u_mem/memory[107] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1215_  (.RESET_B(net93),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0115_ ),
    .Q(\u_ppwm/u_mem/_0000_ ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1216_  (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net296),
    .Q(\u_ppwm/u_mem/_0001_ ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1217_  (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0117_ ),
    .Q(\u_ppwm/u_mem/_0002_ ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1218_  (.RESET_B(net164),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0118_ ),
    .Q(\u_ppwm/u_mem/_0003_ ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1219_  (.RESET_B(net148),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0119_ ),
    .Q(\u_ppwm/u_mem/bit_count[0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1220_  (.RESET_B(net117),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0120_ ),
    .Q(\u_ppwm/u_mem/bit_count[1] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1221_  (.RESET_B(net85),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net613),
    .Q(\u_ppwm/u_mem/bit_count[2] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1222_  (.RESET_B(net172),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0122_ ),
    .Q(\u_ppwm/u_mem/bit_count[3] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1223_  (.RESET_B(net133),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0123_ ),
    .Q(\u_ppwm/u_mem/bit_count[4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1224_  (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net589),
    .Q(\u_ppwm/u_mem/bit_count[5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1225_  (.RESET_B(net175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net567),
    .Q(\u_ppwm/u_mem/bit_count[6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1226_  (.RESET_B(net176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net334),
    .Q(\u_ppwm/u_mem/state_q[0] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1227_  (.RESET_B(net156),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net626),
    .Q(\u_ppwm/mem_write_done ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1228_  (.RESET_B(net101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_mem/_0006_ ),
    .Q(\u_ppwm/u_mem/state_q[2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_tiehi \u_ppwm/u_mem/_1153__56  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net56));
 sg13g2_tiehi \u_ppwm/u_mem/_1208__57  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net57));
 sg13g2_tiehi \u_ppwm/u_mem/_1152__58  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net58));
 sg13g2_tiehi \u_ppwm/u_mem/_1189__59  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net59));
 sg13g2_tiehi \u_ppwm/u_mem/_1151__60  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net60));
 sg13g2_tiehi \u_ppwm/u_mem/_1217__61  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net61));
 sg13g2_tiehi \u_ppwm/u_mem/_1150__62  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net62));
 sg13g2_tiehi \u_ppwm/u_mem/_1188__63  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net63));
 sg13g2_tiehi \u_ppwm/u_mem/_1149__64  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net64));
 sg13g2_tiehi \u_ppwm/u_mem/_1207__65  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net65));
 sg13g2_tiehi \u_ppwm/u_mem/_1148__66  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net66));
 sg13g2_tiehi \u_ppwm/u_mem/_1187__67  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net67));
 sg13g2_tiehi \u_ppwm/u_mem/_1147__68  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net68));
 sg13g2_tiehi \u_ppwm/u_mem/_1224__69  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net69));
 sg13g2_tiehi \u_ppwm/u_mem/_1146__70  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net70));
 sg13g2_tiehi \u_ppwm/u_mem/_1186__71  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net71));
 sg13g2_tiehi \u_ppwm/u_mem/_1145__72  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net72));
 sg13g2_tiehi \u_ppwm/u_mem/_1206__73  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net73));
 sg13g2_tiehi \u_ppwm/u_mem/_1144__74  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net74));
 sg13g2_tiehi \u_ppwm/u_mem/_1185__75  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net75));
 sg13g2_tiehi \u_ppwm/u_mem/_1143__76  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net76));
 sg13g2_tiehi \u_ppwm/u_mem/_1216__77  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net77));
 sg13g2_tiehi \u_ppwm/u_mem/_1142__78  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net78));
 sg13g2_tiehi \u_ppwm/u_mem/_1184__79  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net79));
 sg13g2_tiehi \u_ppwm/u_mem/_1141__80  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net80));
 sg13g2_tiehi \u_ppwm/u_mem/_1205__81  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net81));
 sg13g2_tiehi \u_ppwm/u_mem/_1140__82  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net82));
 sg13g2_tiehi \u_ppwm/u_mem/_1183__83  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net83));
 sg13g2_tiehi \u_ppwm/u_mem/_1139__84  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net84));
 sg13g2_tiehi \u_ppwm/u_mem/_1221__85  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net85));
 sg13g2_tiehi \u_ppwm/u_mem/_1138__86  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net86));
 sg13g2_tiehi \u_ppwm/u_mem/_1182__87  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net87));
 sg13g2_tiehi \u_ppwm/u_mem/_1137__88  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net88));
 sg13g2_tiehi \u_ppwm/u_mem/_1204__89  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net89));
 sg13g2_tiehi \u_ppwm/u_mem/_1136__90  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net90));
 sg13g2_tiehi \u_ppwm/u_mem/_1181__91  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net91));
 sg13g2_tiehi \u_ppwm/u_mem/_1135__92  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net92));
 sg13g2_tiehi \u_ppwm/u_mem/_1215__93  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net93));
 sg13g2_tiehi \u_ppwm/u_mem/_1134__94  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net94));
 sg13g2_tiehi \u_ppwm/u_mem/_1180__95  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net95));
 sg13g2_tiehi \u_ppwm/u_mem/_1133__96  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net96));
 sg13g2_tiehi \u_ppwm/u_mem/_1203__97  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net97));
 sg13g2_tiehi \u_ppwm/u_mem/_1132__98  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net98));
 sg13g2_tiehi \u_ppwm/u_mem/_1179__99  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net99));
 sg13g2_tiehi \u_ppwm/u_mem/_1131__100  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net100));
 sg13g2_tiehi \u_ppwm/u_mem/_1228__101  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net101));
 sg13g2_tiehi \u_ppwm/u_mem/_1130__102  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net102));
 sg13g2_tiehi \u_ppwm/u_mem/_1178__103  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net103));
 sg13g2_tiehi \u_ppwm/u_mem/_1129__104  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net104));
 sg13g2_tiehi \u_ppwm/u_mem/_1202__105  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net105));
 sg13g2_tiehi \u_ppwm/u_mem/_1128__106  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net106));
 sg13g2_tiehi \u_ppwm/u_mem/_1177__107  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net107));
 sg13g2_tiehi \u_ppwm/u_mem/_1127__108  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net108));
 sg13g2_tiehi \u_ppwm/u_mem/_1214__109  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net109));
 sg13g2_tiehi \u_ppwm/u_mem/_1126__110  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net110));
 sg13g2_tiehi \u_ppwm/u_mem/_1176__111  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net111));
 sg13g2_tiehi \u_ppwm/u_mem/_1125__112  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net112));
 sg13g2_tiehi \u_ppwm/u_mem/_1201__113  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net113));
 sg13g2_tiehi \u_ppwm/u_mem/_1124__114  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net114));
 sg13g2_tiehi \u_ppwm/u_mem/_1175__115  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net115));
 sg13g2_tiehi \u_ppwm/u_mem/_1123__116  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net116));
 sg13g2_tiehi \u_ppwm/u_mem/_1220__117  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net117));
 sg13g2_tiehi \u_ppwm/u_mem/_1122__118  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net118));
 sg13g2_tiehi \u_ppwm/u_mem/_1174__119  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net119));
 sg13g2_tiehi \u_ppwm/u_mem/_1121__120  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net120));
 sg13g2_tiehi \u_ppwm/u_mem/_1200__121  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net121));
 sg13g2_tiehi \u_ppwm/u_mem/_1120__122  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net122));
 sg13g2_tiehi \u_ppwm/u_mem/_1173__123  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net123));
 sg13g2_tiehi \u_ppwm/u_mem/_1119__124  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net124));
 sg13g2_tiehi \u_ppwm/u_mem/_1213__125  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net125));
 sg13g2_tiehi \u_ppwm/u_mem/_1118__126  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net126));
 sg13g2_tiehi \u_ppwm/u_mem/_1172__127  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net127));
 sg13g2_tiehi \u_ppwm/u_mem/_1117__128  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net128));
 sg13g2_tiehi \u_ppwm/u_mem/_1199__129  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net129));
 sg13g2_tiehi \u_ppwm/u_mem/_1116__130  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net130));
 sg13g2_tiehi \u_ppwm/u_mem/_1171__131  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net131));
 sg13g2_tiehi \u_ppwm/u_mem/_1115__132  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net132));
 sg13g2_tiehi \u_ppwm/u_mem/_1223__133  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net133));
 sg13g2_tiehi \u_ppwm/u_mem/_1114__134  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net134));
 sg13g2_tiehi \u_ppwm/u_mem/_1170__135  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net135));
 sg13g2_tiehi \u_ppwm/u_mem/_1113__136  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net136));
 sg13g2_tiehi \u_ppwm/u_mem/_1198__137  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net137));
 sg13g2_tiehi \u_ppwm/u_mem/_1112__138  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net138));
 sg13g2_tiehi \u_ppwm/u_mem/_1169__139  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net139));
 sg13g2_tiehi \u_ppwm/u_mem/_1111__140  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net140));
 sg13g2_tiehi \u_ppwm/u_mem/_1212__141  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net141));
 sg13g2_tiehi \u_ppwm/u_mem/_1110__142  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net142));
 sg13g2_tiehi \u_ppwm/u_mem/_1168__143  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net143));
 sg13g2_tiehi \u_ppwm/u_mem/_1109__144  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net144));
 sg13g2_tiehi \u_ppwm/u_mem/_1197__145  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net145));
 sg13g2_tiehi \u_ppwm/u_mem/_1108__146  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net146));
 sg13g2_tiehi \u_ppwm/u_mem/_1167__147  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net147));
 sg13g2_tiehi \u_ppwm/u_mem/_1219__148  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net148));
 sg13g2_tiehi \u_ppwm/u_mem/_1166__149  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net149));
 sg13g2_tiehi \u_ppwm/u_mem/_1196__150  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net150));
 sg13g2_tiehi \u_ppwm/u_mem/_1165__151  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net151));
 sg13g2_tiehi \u_ppwm/u_mem/_1211__152  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net152));
 sg13g2_tiehi \u_ppwm/u_mem/_1164__153  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net153));
 sg13g2_tiehi \u_ppwm/u_mem/_1195__154  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net154));
 sg13g2_tiehi \u_ppwm/u_mem/_1163__155  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net155));
 sg13g2_tiehi \u_ppwm/u_mem/_1227__156  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net156));
 sg13g2_tiehi \u_ppwm/u_mem/_1162__157  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net157));
 sg13g2_tiehi \u_ppwm/u_mem/_1194__158  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net158));
 sg13g2_tiehi \u_ppwm/u_mem/_1161__159  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net159));
 sg13g2_tiehi \u_ppwm/u_mem/_1210__160  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net160));
 sg13g2_tiehi \u_ppwm/u_mem/_1160__161  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net161));
 sg13g2_tiehi \u_ppwm/u_mem/_1193__162  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net162));
 sg13g2_tiehi \u_ppwm/u_mem/_1159__163  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net163));
 sg13g2_tiehi \u_ppwm/u_mem/_1218__164  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net164));
 sg13g2_tiehi \u_ppwm/u_mem/_1158__165  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net165));
 sg13g2_tiehi \u_ppwm/u_mem/_1192__166  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net166));
 sg13g2_tiehi \u_ppwm/u_mem/_1157__167  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net167));
 sg13g2_tiehi \u_ppwm/u_mem/_1209__168  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net168));
 sg13g2_tiehi \u_ppwm/u_mem/_1156__169  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net169));
 sg13g2_tiehi \u_ppwm/u_mem/_1191__170  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net170));
 sg13g2_tiehi \u_ppwm/u_mem/_1155__171  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net171));
 sg13g2_tiehi \u_ppwm/u_mem/_1222__172  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net172));
 sg13g2_tiehi \u_ppwm/u_mem/_1154__173  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net173));
 sg13g2_tiehi \u_ppwm/u_mem/_1107__174  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net174));
 sg13g2_tiehi \u_ppwm/u_mem/_1225__175  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net175));
 sg13g2_tiehi \u_ppwm/u_mem/_1226__176  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net176));
 sg13g2_tiehi \u_ppwm/u_pwm/_234__177  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net177));
 sg13g2_inv_1 \u_ppwm/u_pwm/_125_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_072_ ),
    .A(net593),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_126_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_073_ ),
    .A(net299),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_127_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_074_ ),
    .A(net238),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_128_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_075_ ),
    .A(net211),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_129_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_076_ ),
    .A(net209),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_130_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_077_ ),
    .A(net260),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_pwm/_131_  (.Y(\u_ppwm/u_pwm/_078_ ),
    .A(net207),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_132_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_079_ ),
    .A(net533),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_133_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_080_ ),
    .A(net203),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_134_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_081_ ),
    .A(net215),
    .VSS(VGND));
 sg13g2_inv_1 \u_ppwm/u_pwm/_135_  (.VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_082_ ),
    .A(net199),
    .VSS(VGND));
 sg13g2_inv_2 \u_ppwm/u_pwm/_136_  (.Y(\u_ppwm/u_pwm/_083_ ),
    .A(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 \u_ppwm/u_pwm/_137_  (.A(\u_ppwm/u_pwm/counter[3] ),
    .B(\u_ppwm/u_pwm/counter[2] ),
    .C(\u_ppwm/u_pwm/counter[1] ),
    .D(\u_ppwm/u_pwm/counter[0] ),
    .Y(\u_ppwm/u_pwm/_084_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_138_  (.A(\u_ppwm/u_pwm/counter[9] ),
    .B(\u_ppwm/u_pwm/counter[8] ),
    .Y(\u_ppwm/u_pwm/_085_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 \u_ppwm/u_pwm/_139_  (.A(\u_ppwm/u_pwm/counter[7] ),
    .B(\u_ppwm/u_pwm/counter[6] ),
    .C(\u_ppwm/u_pwm/counter[5] ),
    .D(\u_ppwm/u_pwm/counter[4] ),
    .Y(\u_ppwm/u_pwm/_086_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_pwm/_140_  (.B(\u_ppwm/u_pwm/_085_ ),
    .C(\u_ppwm/u_pwm/_086_ ),
    .A(\u_ppwm/u_pwm/_084_ ),
    .Y(\u_ppwm/u_pwm/_087_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_141_  (.B1(net492),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_088_ ),
    .VSS(VGND),
    .A1(net466),
    .A2(net390));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_142_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_082_ ),
    .A2(net390),
    .Y(\u_ppwm/u_pwm/_000_ ),
    .B1(\u_ppwm/u_pwm/_088_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_143_  (.B1(net492),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_089_ ),
    .VSS(VGND),
    .A1(net465),
    .A2(net390));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_144_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_081_ ),
    .A2(net390),
    .Y(\u_ppwm/u_pwm/_001_ ),
    .B1(\u_ppwm/u_pwm/_089_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_145_  (.B1(net493),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_090_ ),
    .VSS(VGND),
    .A1(net463),
    .A2(net390));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_146_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_080_ ),
    .A2(net391),
    .Y(\u_ppwm/u_pwm/_002_ ),
    .B1(\u_ppwm/u_pwm/_090_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_147_  (.B1(net490),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_091_ ),
    .VSS(VGND),
    .A1(\u_ppwm/pwm_value[3] ),
    .A2(net390));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_148_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_079_ ),
    .A2(net390),
    .Y(\u_ppwm/u_pwm/_003_ ),
    .B1(\u_ppwm/u_pwm/_091_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_149_  (.B1(net490),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_092_ ),
    .VSS(VGND),
    .A1(net460),
    .A2(net389));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_150_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_078_ ),
    .A2(net389),
    .Y(\u_ppwm/u_pwm/_004_ ),
    .B1(\u_ppwm/u_pwm/_092_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_151_  (.B1(net490),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_093_ ),
    .VSS(VGND),
    .A1(net458),
    .A2(net389));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_152_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_077_ ),
    .A2(net389),
    .Y(\u_ppwm/u_pwm/_005_ ),
    .B1(\u_ppwm/u_pwm/_093_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_153_  (.B1(net490),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_094_ ),
    .VSS(VGND),
    .A1(net456),
    .A2(net389));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_154_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_076_ ),
    .A2(net391),
    .Y(\u_ppwm/u_pwm/_006_ ),
    .B1(\u_ppwm/u_pwm/_094_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_155_  (.B1(net490),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_095_ ),
    .VSS(VGND),
    .A1(\u_ppwm/pwm_value[7] ),
    .A2(net389));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_156_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_075_ ),
    .A2(net391),
    .Y(\u_ppwm/u_pwm/_007_ ),
    .B1(\u_ppwm/u_pwm/_095_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_157_  (.B1(net490),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_096_ ),
    .VSS(VGND),
    .A1(net455),
    .A2(net389));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_158_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_074_ ),
    .A2(net389),
    .Y(\u_ppwm/u_pwm/_008_ ),
    .B1(\u_ppwm/u_pwm/_096_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_159_  (.B1(net490),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_097_ ),
    .VSS(VGND),
    .A1(net454),
    .A2(net391));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_160_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_073_ ),
    .A2(net390),
    .Y(\u_ppwm/u_pwm/_009_ ),
    .B1(\u_ppwm/u_pwm/_097_ ));
 sg13g2_and2_1 \u_ppwm/u_pwm/_161_  (.A(net625),
    .B(net647),
    .X(\u_ppwm/u_pwm/_098_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_162_  (.B1(net489),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_099_ ),
    .VSS(VGND),
    .A1(net625),
    .A2(net647));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_163_  (.A(\u_ppwm/u_pwm/_098_ ),
    .B(\u_ppwm/u_pwm/_099_ ),
    .Y(\u_ppwm/u_pwm/_010_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_164_  (.B1(net489),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_100_ ),
    .VSS(VGND),
    .A1(net549),
    .A2(\u_ppwm/u_pwm/_098_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_165_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net549),
    .A2(\u_ppwm/u_pwm/_098_ ),
    .Y(\u_ppwm/u_pwm/_011_ ),
    .B1(\u_ppwm/u_pwm/_100_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_166_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(net549),
    .A2(\u_ppwm/u_pwm/_098_ ),
    .Y(\u_ppwm/u_pwm/_101_ ),
    .B1(net572));
 sg13g2_and4_1 \u_ppwm/u_pwm/_167_  (.A(net625),
    .B(net572),
    .C(net549),
    .D(net647),
    .X(\u_ppwm/u_pwm/_102_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_pwm/_168_  (.A(\u_ppwm/u_pwm/_083_ ),
    .B(net573),
    .C(\u_ppwm/u_pwm/_102_ ),
    .Y(\u_ppwm/u_pwm/_012_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_169_  (.A(net651),
    .B(\u_ppwm/u_pwm/_102_ ),
    .Y(\u_ppwm/u_pwm/_022_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 \u_ppwm/u_pwm/_170_  (.A(net651),
    .B(\u_ppwm/u_pwm/_102_ ),
    .X(\u_ppwm/u_pwm/_023_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_pwm/_171_  (.A(\u_ppwm/u_pwm/_083_ ),
    .B(\u_ppwm/u_pwm/_022_ ),
    .C(\u_ppwm/u_pwm/_023_ ),
    .Y(\u_ppwm/u_pwm/_013_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_pwm/_172_  (.Y(\u_ppwm/u_pwm/_024_ ),
    .A(net652),
    .B(\u_ppwm/u_pwm/_023_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_173_  (.A(\u_ppwm/u_pwm/_083_ ),
    .B(\u_ppwm/u_pwm/_024_ ),
    .Y(\u_ppwm/u_pwm/_014_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_174_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/counter[4] ),
    .A2(\u_ppwm/u_pwm/_023_ ),
    .Y(\u_ppwm/u_pwm/_025_ ),
    .B1(net601));
 sg13g2_and3_2 \u_ppwm/u_pwm/_175_  (.X(\u_ppwm/u_pwm/_026_ ),
    .A(net601),
    .B(net652),
    .C(\u_ppwm/u_pwm/_023_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_pwm/_176_  (.A(\u_ppwm/u_pwm/_083_ ),
    .B(net602),
    .C(\u_ppwm/u_pwm/_026_ ),
    .Y(\u_ppwm/u_pwm/_015_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \u_ppwm/u_pwm/_177_  (.Y(\u_ppwm/u_pwm/_027_ ),
    .A(net636),
    .B(\u_ppwm/u_pwm/_026_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_178_  (.A(\u_ppwm/u_pwm/_083_ ),
    .B(\u_ppwm/u_pwm/_027_ ),
    .Y(\u_ppwm/u_pwm/_016_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_179_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/counter[6] ),
    .A2(\u_ppwm/u_pwm/_026_ ),
    .Y(\u_ppwm/u_pwm/_028_ ),
    .B1(net546));
 sg13g2_nand3_1 \u_ppwm/u_pwm/_180_  (.B(net636),
    .C(\u_ppwm/u_pwm/_026_ ),
    .A(net546),
    .Y(\u_ppwm/u_pwm/_029_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_181_  (.Y(\u_ppwm/u_pwm/_030_ ),
    .A(net489),
    .B(\u_ppwm/u_pwm/_029_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_182_  (.A(net547),
    .B(\u_ppwm/u_pwm/_030_ ),
    .Y(\u_ppwm/u_pwm/_017_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 \u_ppwm/u_pwm/_183_  (.VSS(VGND),
    .VDD(VPWR),
    .X(\u_ppwm/u_pwm/_031_ ),
    .B(\u_ppwm/u_pwm/_029_ ),
    .A(\u_ppwm/u_pwm/_072_ ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_184_  (.Y(\u_ppwm/u_pwm/_032_ ),
    .A(net489),
    .B(\u_ppwm/u_pwm/_031_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_185_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_072_ ),
    .A2(net637),
    .Y(\u_ppwm/u_pwm/_018_ ),
    .B1(\u_ppwm/u_pwm/_032_ ));
 sg13g2_nand4_1 \u_ppwm/u_pwm/_186_  (.B(net593),
    .C(net546),
    .A(\u_ppwm/u_pwm/counter[9] ),
    .Y(\u_ppwm/u_pwm/_033_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_pwm/counter[6] ));
 sg13g2_xor2_1 \u_ppwm/u_pwm/_187_  (.B(\u_ppwm/u_pwm/_031_ ),
    .A(net644),
    .X(\u_ppwm/u_pwm/_034_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_188_  (.A(\u_ppwm/u_pwm/_083_ ),
    .B(\u_ppwm/u_pwm/_034_ ),
    .Y(\u_ppwm/u_pwm/_019_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 \u_ppwm/u_pwm/_189_  (.B(\u_ppwm/u_pwm/counter[0] ),
    .C(net489),
    .A(net549),
    .Y(\u_ppwm/u_pwm/_035_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_pwm/_190_  (.B(\u_ppwm/u_pwm/counter[4] ),
    .C(\u_ppwm/u_pwm/counter[3] ),
    .A(\u_ppwm/u_pwm/counter[5] ),
    .Y(\u_ppwm/u_pwm/_036_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net572));
 sg13g2_nor3_1 \u_ppwm/u_pwm/_191_  (.A(net594),
    .B(\u_ppwm/u_pwm/_035_ ),
    .C(\u_ppwm/u_pwm/_036_ ),
    .Y(\u_ppwm/u_pwm/_020_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_192_  (.A(\u_ppwm/u_pwm/cmp_value[2] ),
    .B_N(\u_ppwm/u_pwm/counter[2] ),
    .Y(\u_ppwm/u_pwm/_037_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_193_  (.A(\u_ppwm/u_pwm/cmp_value[3] ),
    .B_N(\u_ppwm/u_pwm/counter[3] ),
    .Y(\u_ppwm/u_pwm/_038_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_194_  (.A(\u_ppwm/u_pwm/counter[3] ),
    .B_N(\u_ppwm/u_pwm/cmp_value[3] ),
    .Y(\u_ppwm/u_pwm/_039_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_195_  (.Y(\u_ppwm/u_pwm/_040_ ),
    .B(\u_ppwm/u_pwm/cmp_value[3] ),
    .A_N(\u_ppwm/u_pwm/counter[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_196_  (.B1(\u_ppwm/u_pwm/_040_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_041_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_pwm/_037_ ),
    .A2(\u_ppwm/u_pwm/_038_ ));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_197_  (.A(\u_ppwm/u_pwm/cmp_value[1] ),
    .B_N(\u_ppwm/u_pwm/counter[1] ),
    .Y(\u_ppwm/u_pwm/_042_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_198_  (.Y(\u_ppwm/u_pwm/_043_ ),
    .B(\u_ppwm/u_pwm/cmp_value[0] ),
    .A_N(\u_ppwm/u_pwm/counter[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_199_  (.Y(\u_ppwm/u_pwm/_044_ ),
    .B(\u_ppwm/u_pwm/cmp_value[1] ),
    .A_N(\u_ppwm/u_pwm/counter[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_200_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_043_ ),
    .A2(\u_ppwm/u_pwm/_044_ ),
    .Y(\u_ppwm/u_pwm/_045_ ),
    .B1(\u_ppwm/u_pwm/_042_ ));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_201_  (.A(\u_ppwm/u_pwm/counter[2] ),
    .B_N(\u_ppwm/u_pwm/cmp_value[2] ),
    .Y(\u_ppwm/u_pwm/_046_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 \u_ppwm/u_pwm/_202_  (.A(\u_ppwm/u_pwm/_037_ ),
    .B(\u_ppwm/u_pwm/_038_ ),
    .C(\u_ppwm/u_pwm/_039_ ),
    .D(\u_ppwm/u_pwm/_046_ ),
    .X(\u_ppwm/u_pwm/_047_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_203_  (.B1(\u_ppwm/u_pwm/_041_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_048_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_pwm/_045_ ),
    .A2(\u_ppwm/u_pwm/_047_ ));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_204_  (.Y(\u_ppwm/u_pwm/_049_ ),
    .B(\u_ppwm/u_pwm/counter[7] ),
    .A_N(\u_ppwm/u_pwm/cmp_value[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_205_  (.Y(\u_ppwm/u_pwm/_050_ ),
    .B(\u_ppwm/u_pwm/counter[6] ),
    .A_N(\u_ppwm/u_pwm/cmp_value[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_206_  (.Y(\u_ppwm/u_pwm/_051_ ),
    .A(\u_ppwm/u_pwm/_049_ ),
    .B(\u_ppwm/u_pwm/_050_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_207_  (.Y(\u_ppwm/u_pwm/_052_ ),
    .B(\u_ppwm/u_pwm/cmp_value[6] ),
    .A_N(\u_ppwm/u_pwm/counter[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_208_  (.Y(\u_ppwm/u_pwm/_053_ ),
    .B(\u_ppwm/u_pwm/cmp_value[7] ),
    .A_N(\u_ppwm/u_pwm/counter[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 \u_ppwm/u_pwm/_209_  (.B(\u_ppwm/u_pwm/_050_ ),
    .C(\u_ppwm/u_pwm/_052_ ),
    .A(\u_ppwm/u_pwm/_049_ ),
    .Y(\u_ppwm/u_pwm/_054_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_ppwm/u_pwm/_053_ ));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_210_  (.A(\u_ppwm/u_pwm/cmp_value[5] ),
    .B_N(\u_ppwm/u_pwm/counter[5] ),
    .Y(\u_ppwm/u_pwm/_055_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_211_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/counter[4] ),
    .A2(\u_ppwm/u_pwm/_078_ ),
    .Y(\u_ppwm/u_pwm/_056_ ),
    .B1(\u_ppwm/u_pwm/_055_ ));
 sg13g2_a21o_1 \u_ppwm/u_pwm/_212_  (.A2(\u_ppwm/u_pwm/_078_ ),
    .A1(\u_ppwm/u_pwm/counter[4] ),
    .B1(\u_ppwm/u_pwm/_055_ ),
    .X(\u_ppwm/u_pwm/_057_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_213_  (.A(\u_ppwm/u_pwm/counter[4] ),
    .B(\u_ppwm/u_pwm/_078_ ),
    .Y(\u_ppwm/u_pwm/_058_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_214_  (.A(\u_ppwm/u_pwm/counter[5] ),
    .B(\u_ppwm/u_pwm/_077_ ),
    .Y(\u_ppwm/u_pwm/_059_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 \u_ppwm/u_pwm/_215_  (.A(\u_ppwm/u_pwm/_054_ ),
    .B(\u_ppwm/u_pwm/_057_ ),
    .C(\u_ppwm/u_pwm/_058_ ),
    .D(\u_ppwm/u_pwm/_059_ ),
    .Y(\u_ppwm/u_pwm/_060_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 \u_ppwm/u_pwm/_216_  (.A(\u_ppwm/u_pwm/_054_ ),
    .B(\u_ppwm/u_pwm/_056_ ),
    .C(\u_ppwm/u_pwm/_059_ ),
    .Y(\u_ppwm/u_pwm/_061_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 \u_ppwm/u_pwm/_217_  (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_ppwm/u_pwm/_048_ ),
    .C1(\u_ppwm/u_pwm/_061_ ),
    .B1(\u_ppwm/u_pwm/_060_ ),
    .A1(\u_ppwm/u_pwm/_051_ ),
    .Y(\u_ppwm/u_pwm/_062_ ),
    .A2(\u_ppwm/u_pwm/_053_ ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_218_  (.Y(\u_ppwm/u_pwm/_063_ ),
    .A(\u_ppwm/u_pwm/counter[8] ),
    .B(\u_ppwm/u_pwm/_074_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_219_  (.A(net644),
    .B(\u_ppwm/u_pwm/_073_ ),
    .Y(\u_ppwm/u_pwm/_064_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_220_  (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_ppwm/u_pwm/_072_ ),
    .A2(\u_ppwm/u_pwm/cmp_value[8] ),
    .Y(\u_ppwm/u_pwm/_065_ ),
    .B1(\u_ppwm/u_pwm/_064_ ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_221_  (.Y(\u_ppwm/u_pwm/_066_ ),
    .A(\u_ppwm/u_pwm/_063_ ),
    .B(\u_ppwm/u_pwm/_065_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_222_  (.A(\u_ppwm/u_pwm/_062_ ),
    .B(\u_ppwm/u_pwm/_066_ ),
    .Y(\u_ppwm/u_pwm/_067_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_223_  (.Y(\u_ppwm/u_pwm/_068_ ),
    .A(net644),
    .B(\u_ppwm/u_pwm/_073_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_224_  (.B1(\u_ppwm/u_pwm/_068_ ),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_069_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_pwm/_063_ ),
    .A2(\u_ppwm/u_pwm/_064_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_225_  (.B1(net247),
    .VDD(VPWR),
    .Y(\u_ppwm/u_pwm/_070_ ),
    .VSS(VGND),
    .A1(\u_ppwm/u_pwm/_067_ ),
    .A2(\u_ppwm/u_pwm/_069_ ));
 sg13g2_or3_1 \u_ppwm/u_pwm/_226_  (.A(net247),
    .B(\u_ppwm/u_pwm/_067_ ),
    .C(\u_ppwm/u_pwm/_069_ ),
    .X(\u_ppwm/u_pwm/_071_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 \u_ppwm/u_pwm/_227_  (.X(\u_ppwm/u_pwm/_021_ ),
    .A(net489),
    .B(\u_ppwm/u_pwm/_070_ ),
    .C(\u_ppwm/u_pwm/_071_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_228_  (.RESET_B(net190),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net200),
    .Q(\u_ppwm/u_pwm/cmp_value[0] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_229_  (.RESET_B(net187),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net216),
    .Q(\u_ppwm/u_pwm/cmp_value[1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_230_  (.RESET_B(net185),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net204),
    .Q(\u_ppwm/u_pwm/cmp_value[2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_231_  (.RESET_B(net183),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net534),
    .Q(\u_ppwm/u_pwm/cmp_value[3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_232_  (.RESET_B(net181),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net208),
    .Q(\u_ppwm/u_pwm/cmp_value[4] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_233_  (.RESET_B(net179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net261),
    .Q(\u_ppwm/u_pwm/cmp_value[5] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_234_  (.RESET_B(net177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net210),
    .Q(\u_ppwm/u_pwm/cmp_value[6] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_235_  (.RESET_B(net197),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net212),
    .Q(\u_ppwm/u_pwm/cmp_value[7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_236_  (.RESET_B(net195),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net239),
    .Q(\u_ppwm/u_pwm/cmp_value[8] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_237_  (.RESET_B(net193),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net300),
    .Q(\u_ppwm/u_pwm/cmp_value[9] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_238_  (.RESET_B(net191),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_pwm/_010_ ),
    .Q(\u_ppwm/u_pwm/counter[0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_239_  (.RESET_B(net189),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net550),
    .Q(\u_ppwm/u_pwm/counter[1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_240_  (.RESET_B(net186),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net574),
    .Q(\u_ppwm/u_pwm/counter[2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_241_  (.RESET_B(net182),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_pwm/_013_ ),
    .Q(\u_ppwm/u_pwm/counter[3] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_242_  (.RESET_B(net178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_pwm/_014_ ),
    .Q(\u_ppwm/u_pwm/counter[4] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_243_  (.RESET_B(net196),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net603),
    .Q(\u_ppwm/u_pwm/counter[5] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_244_  (.RESET_B(net192),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_pwm/_016_ ),
    .Q(\u_ppwm/u_pwm/counter[6] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_245_  (.RESET_B(net188),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net548),
    .Q(\u_ppwm/u_pwm/counter[7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_246_  (.RESET_B(net180),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_pwm/_018_ ),
    .Q(\u_ppwm/u_pwm/counter[8] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_247_  (.RESET_B(net194),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_pwm/_019_ ),
    .Q(\u_ppwm/u_pwm/counter[9] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_248_  (.RESET_B(net184),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net595),
    .Q(\u_ppwm/period_start ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_249_  (.RESET_B(net198),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\u_ppwm/u_pwm/_021_ ),
    .Q(net2),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_tiehi \u_ppwm/u_pwm/_242__178  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net178));
 sg13g2_tiehi \u_ppwm/u_pwm/_233__179  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net179));
 sg13g2_tiehi \u_ppwm/u_pwm/_246__180  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net180));
 sg13g2_tiehi \u_ppwm/u_pwm/_232__181  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net181));
 sg13g2_tiehi \u_ppwm/u_pwm/_241__182  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net182));
 sg13g2_tiehi \u_ppwm/u_pwm/_231__183  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net183));
 sg13g2_tiehi \u_ppwm/u_pwm/_248__184  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net184));
 sg13g2_tiehi \u_ppwm/u_pwm/_230__185  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net185));
 sg13g2_tiehi \u_ppwm/u_pwm/_240__186  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net186));
 sg13g2_tiehi \u_ppwm/u_pwm/_229__187  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net187));
 sg13g2_tiehi \u_ppwm/u_pwm/_245__188  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net188));
 sg13g2_tiehi \u_ppwm/u_pwm/_239__189  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net189));
 sg13g2_tiehi \u_ppwm/u_pwm/_228__190  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net190));
 sg13g2_tiehi \u_ppwm/u_pwm/_238__191  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net191));
 sg13g2_tiehi \u_ppwm/u_pwm/_244__192  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net192));
 sg13g2_tiehi \u_ppwm/u_pwm/_237__193  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net193));
 sg13g2_tiehi \u_ppwm/u_pwm/_247__194  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net194));
 sg13g2_tiehi \u_ppwm/u_pwm/_236__195  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net195));
 sg13g2_tiehi \u_ppwm/u_pwm/_243__196  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net196));
 sg13g2_tiehi \u_ppwm/u_pwm/_235__197  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net197));
 sg13g2_tiehi \u_ppwm/u_pwm/_249__198  (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net198));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout349 (.A(net351),
    .X(net349),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout350 (.A(net351),
    .X(net350),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout351 (.A(\u_ppwm/u_ex/_0419_ ),
    .X(net351),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout352 (.A(net353),
    .X(net352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout353 (.A(net354),
    .X(net353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout354 (.A(\u_ppwm/u_ex/_0251_ ),
    .X(net354),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout355 (.A(\u_ppwm/u_ex/_0413_ ),
    .X(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout356 (.A(\u_ppwm/u_ex/_0188_ ),
    .X(net356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout357 (.A(net358),
    .X(net357),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout358 (.A(\u_ppwm/u_ex/_0225_ ),
    .X(net358),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout359 (.A(\u_ppwm/u_ex/_0220_ ),
    .X(net359),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout360 (.A(\u_ppwm/u_ex/_0220_ ),
    .X(net360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout361 (.A(\u_ppwm/u_ex/_0220_ ),
    .X(net361),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout362 (.A(net363),
    .X(net362),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout363 (.A(\u_ppwm/u_ex/_0187_ ),
    .X(net363),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout364 (.A(\u_ppwm/u_ex/_0161_ ),
    .X(net364),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout365 (.A(\u_ppwm/u_ex/_0161_ ),
    .X(net365),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout366 (.A(\u_ppwm/u_ex/_0136_ ),
    .X(net366),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout367 (.A(\u_ppwm/u_ex/_0136_ ),
    .X(net367),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout368 (.A(net369),
    .X(net368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout369 (.A(\u_ppwm/u_ex/_0051_ ),
    .X(net369),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout370 (.A(\u_ppwm/u_ex/_0036_ ),
    .X(net370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout371 (.A(net372),
    .X(net371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout372 (.A(net374),
    .X(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout373 (.A(net374),
    .X(net373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout374 (.A(\u_ppwm/instr[6] ),
    .X(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout375 (.A(\u_ppwm/instr[6] ),
    .X(net375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout376 (.A(\u_ppwm/instr[6] ),
    .X(net376),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout377 (.A(net378),
    .X(net377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout378 (.A(net379),
    .X(net378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout379 (.A(net380),
    .X(net379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout380 (.A(\u_ppwm/instr[5] ),
    .X(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout381 (.A(net383),
    .X(net381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout382 (.A(net383),
    .X(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout383 (.A(\u_ppwm/instr[4] ),
    .X(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout384 (.A(net385),
    .X(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout385 (.A(net387),
    .X(net385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout386 (.A(net387),
    .X(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout387 (.A(\u_ppwm/instr[3] ),
    .X(net387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout388 (.A(\u_ppwm/instr[2] ),
    .X(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout389 (.A(net391),
    .X(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout390 (.A(net391),
    .X(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout391 (.A(\u_ppwm/u_pwm/_087_ ),
    .X(net391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout392 (.A(\u_ppwm/u_global_counter/_041_ ),
    .X(net392),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout393 (.A(net394),
    .X(net393),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout394 (.A(\u_ppwm/u_mem/_0241_ ),
    .X(net394),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout395 (.A(net396),
    .X(net395),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout396 (.A(net397),
    .X(net396),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout397 (.A(\u_ppwm/u_mem/_0240_ ),
    .X(net397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout398 (.A(net399),
    .X(net398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout399 (.A(net642),
    .X(net399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout400 (.A(net402),
    .X(net400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout401 (.A(net402),
    .X(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout402 (.A(net406),
    .X(net402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout403 (.A(net404),
    .X(net403),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout404 (.A(net405),
    .X(net404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout405 (.A(net406),
    .X(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout406 (.A(net422),
    .X(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout407 (.A(net408),
    .X(net407),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout408 (.A(net422),
    .X(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout409 (.A(net410),
    .X(net409),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout410 (.A(net411),
    .X(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout411 (.A(net422),
    .X(net411),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout412 (.A(net416),
    .X(net412),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout413 (.A(net416),
    .X(net413),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout414 (.A(net415),
    .X(net414),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout415 (.A(net416),
    .X(net415),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout416 (.A(net422),
    .X(net416),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout417 (.A(net418),
    .X(net417),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout418 (.A(net421),
    .X(net418),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout419 (.A(net420),
    .X(net419),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout420 (.A(net421),
    .X(net420),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout421 (.A(net422),
    .X(net421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout422 (.A(\u_ppwm/u_mem/state_q[2] ),
    .X(net422),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout423 (.A(net424),
    .X(net423),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout424 (.A(net425),
    .X(net424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout425 (.A(\u_ppwm/u_mem/state_q[2] ),
    .X(net425),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout426 (.A(net438),
    .X(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout427 (.A(net431),
    .X(net427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout428 (.A(net431),
    .X(net428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout429 (.A(net431),
    .X(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout430 (.A(net431),
    .X(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout431 (.A(net438),
    .X(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout432 (.A(net435),
    .X(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout433 (.A(net435),
    .X(net433),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout434 (.A(net435),
    .X(net434),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout435 (.A(net437),
    .X(net435),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout436 (.A(net437),
    .X(net436),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout437 (.A(net438),
    .X(net437),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout438 (.A(\u_ppwm/u_mem/state_q[2] ),
    .X(net438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout439 (.A(net654),
    .X(net439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout440 (.A(net633),
    .X(net440),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout441 (.A(net639),
    .X(net441),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout442 (.A(net201),
    .X(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout443 (.A(net655),
    .X(net443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout444 (.A(net665),
    .X(net444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout445 (.A(net653),
    .X(net445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout446 (.A(net686),
    .X(net446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout447 (.A(net686),
    .X(net447),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout448 (.A(net671),
    .X(net448),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout449 (.A(net682),
    .X(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout450 (.A(net681),
    .X(net450),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout451 (.A(net668),
    .X(net451),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout452 (.A(\u_ppwm/u_ex/reg_value_q[2] ),
    .X(net452),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout453 (.A(net678),
    .X(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout454 (.A(net675),
    .X(net454),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout455 (.A(net672),
    .X(net455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout456 (.A(net677),
    .X(net456),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout457 (.A(\u_ppwm/pwm_value[6] ),
    .X(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout458 (.A(net669),
    .X(net458),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout459 (.A(\u_ppwm/pwm_value[5] ),
    .X(net459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout460 (.A(net676),
    .X(net460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout461 (.A(\u_ppwm/pwm_value[4] ),
    .X(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout462 (.A(net690),
    .X(net462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout463 (.A(net680),
    .X(net463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout464 (.A(net465),
    .X(net464),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout465 (.A(net687),
    .X(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout466 (.A(\u_ppwm/pwm_value[0] ),
    .X(net466),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout467 (.A(\u_ppwm/pc[3] ),
    .X(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout468 (.A(net683),
    .X(net468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout469 (.A(net673),
    .X(net469),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout470 (.A(\u_ppwm/pc[2] ),
    .X(net470),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout471 (.A(net472),
    .X(net471),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout472 (.A(\u_ppwm/pc[1] ),
    .X(net472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout473 (.A(net475),
    .X(net473),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout474 (.A(net475),
    .X(net474),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout475 (.A(net689),
    .X(net475),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout476 (.A(net479),
    .X(net476),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout477 (.A(net479),
    .X(net477),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout478 (.A(net479),
    .X(net478),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout479 (.A(net487),
    .X(net479),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout480 (.A(net487),
    .X(net480),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout481 (.A(net487),
    .X(net481),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout482 (.A(net483),
    .X(net482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout483 (.A(net486),
    .X(net483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout484 (.A(net486),
    .X(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout485 (.A(net486),
    .X(net485),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout486 (.A(net487),
    .X(net486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout487 (.A(\u_ppwm/pc[0] ),
    .X(net487),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout488 (.A(net489),
    .X(net488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout489 (.A(net493),
    .X(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout490 (.A(net492),
    .X(net490),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout491 (.A(net492),
    .X(net491),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout492 (.A(net493),
    .X(net492),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout493 (.A(rst_n),
    .X(net493),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout494 (.A(net495),
    .X(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout495 (.A(net500),
    .X(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout496 (.A(net499),
    .X(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout497 (.A(net499),
    .X(net497),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout498 (.A(net499),
    .X(net498),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout499 (.A(net500),
    .X(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout500 (.A(net504),
    .X(net500),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout501 (.A(net504),
    .X(net501),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout502 (.A(net503),
    .X(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout503 (.A(net504),
    .X(net503),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout504 (.A(rst_n),
    .X(net504),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout505 (.A(net506),
    .X(net505),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout506 (.A(net518),
    .X(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout507 (.A(net509),
    .X(net507),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout508 (.A(net509),
    .X(net508),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout509 (.A(net518),
    .X(net509),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout510 (.A(net511),
    .X(net510),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout511 (.A(net512),
    .X(net511),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout512 (.A(net518),
    .X(net512),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout513 (.A(net517),
    .X(net513),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout514 (.A(net517),
    .X(net514),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout515 (.A(net517),
    .X(net515),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout516 (.A(net517),
    .X(net516),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout517 (.A(net518),
    .X(net517),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout518 (.A(rst_n),
    .X(net518),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_ppwm_3 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net3));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload0 (.VDD(VPWR),
    .A(clknet_5_1__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload1 (.A(clknet_5_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload2 (.A(clknet_5_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload3 (.A(clknet_5_14__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload4 (.A(clknet_5_16__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload5 (.A(clknet_5_18__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload6 (.A(clknet_5_20__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload7 (.A(clknet_5_22__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload8 (.A(clknet_5_24__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload9 (.A(clknet_5_31__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_ppwm/u_pwm/cmp_value[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_ppwm/u_pwm/_000_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_ppwm/global_counter[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold4 (.A(\u_ppwm/u_global_counter/_008_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_ppwm/u_pwm/cmp_value[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_ppwm/u_pwm/_002_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold7 (.A(\u_ppwm/u_mem/memory[91] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold8 (.A(\u_ppwm/u_mem/_0097_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_ppwm/u_pwm/cmp_value[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_ppwm/u_pwm/_004_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_ppwm/u_pwm/cmp_value[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_ppwm/u_pwm/_006_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_ppwm/u_pwm/cmp_value[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_ppwm/u_pwm/_007_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_ppwm/u_mem/memory[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_ppwm/u_mem/_0102_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold17 (.A(\u_ppwm/u_pwm/cmp_value[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_ppwm/u_pwm/_001_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_ppwm/u_ex/state_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold20 (.A(\u_ppwm/u_ex/_0056_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_ppwm/u_ex/_0001_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold22 (.A(\u_ppwm/u_mem/memory[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_ppwm/u_mem/_0042_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_ppwm/u_mem/_0000_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_ppwm/u_mem/_0114_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold26 (.A(\u_ppwm/u_mem/memory[59] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_ppwm/u_mem/_0065_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold28 (.A(\u_ppwm/u_mem/memory[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_ppwm/u_mem/_0039_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold30 (.A(\u_ppwm/u_mem/memory[66] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_ppwm/u_mem/_0072_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold32 (.A(\u_ppwm/u_mem/memory[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_ppwm/u_mem/_0093_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u_ppwm/u_mem/memory[89] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_ppwm/u_mem/_0095_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u_ppwm/u_mem/memory[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_ppwm/u_mem/_0079_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_ppwm/u_mem/memory[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u_ppwm/u_mem/_0086_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold40 (.A(\u_ppwm/u_pwm/cmp_value[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_ppwm/u_pwm/_008_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u_ppwm/u_mem/memory[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_ppwm/u_mem/_0054_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold44 (.A(\u_ppwm/u_mem/memory[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_ppwm/u_mem/_0010_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold46 (.A(\u_ppwm/u_mem/memory[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_ppwm/u_mem/memory[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_ppwm/u_mem/_0057_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_ppwm/polarity ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u_ppwm/u_ex/_0008_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_ppwm/u_mem/memory[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u_ppwm/u_mem/_0085_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_ppwm/u_mem/memory[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u_ppwm/u_mem/_0070_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_ppwm/u_mem/memory[101] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u_ppwm/u_mem/_0107_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u_ppwm/u_mem/memory[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold58 (.A(\u_ppwm/u_mem/_0078_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold59 (.A(\u_ppwm/u_mem/memory[90] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_ppwm/u_mem/memory[100] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold61 (.A(\u_ppwm/u_mem/_0106_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u_ppwm/u_pwm/cmp_value[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold63 (.A(\u_ppwm/u_pwm/_005_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_ppwm/u_mem/memory[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold65 (.A(\u_ppwm/u_mem/_0031_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_ppwm/u_mem/memory[60] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold67 (.A(\u_ppwm/u_mem/memory[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_ppwm/u_mem/_0077_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold69 (.A(\u_ppwm/u_mem/memory[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold70 (.A(\u_ppwm/u_mem/_0069_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold71 (.A(\u_ppwm/u_mem/memory[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold72 (.A(\u_ppwm/u_mem/_0053_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold73 (.A(\u_ppwm/u_mem/memory[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold74 (.A(\u_ppwm/u_mem/_0060_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold75 (.A(\u_ppwm/u_mem/memory[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold76 (.A(\u_ppwm/u_mem/_0046_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold77 (.A(\u_ppwm/u_mem/memory[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_ppwm/u_mem/_0020_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold79 (.A(\u_ppwm/u_mem/memory[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_ppwm/u_mem/memory[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold81 (.A(\u_ppwm/u_mem/_0051_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_ppwm/u_mem/memory[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold83 (.A(\u_ppwm/u_mem/_0017_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_ppwm/u_mem/memory[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold85 (.A(\u_ppwm/u_mem/_0028_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_ppwm/u_mem/memory[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold87 (.A(\u_ppwm/u_mem/_0013_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_ppwm/u_mem/memory[56] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold89 (.A(\u_ppwm/u_mem/_0062_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold90 (.A(\u_ppwm/u_mem/memory[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold91 (.A(\u_ppwm/u_mem/_0034_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_ppwm/u_mem/memory[107] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold93 (.A(\u_ppwm/u_mem/_0113_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold94 (.A(\u_ppwm/u_mem/memory[67] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_ppwm/u_mem/memory[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold96 (.A(\u_ppwm/u_mem/_0019_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_ppwm/u_mem/_0002_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold98 (.A(\u_ppwm/u_mem/_0116_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold99 (.A(\u_ppwm/u_mem/memory[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold100 (.A(\u_ppwm/u_mem/memory[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold101 (.A(\u_ppwm/u_pwm/cmp_value[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_ppwm/u_pwm/_009_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold103 (.A(\u_ppwm/u_mem/memory[99] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold104 (.A(\u_ppwm/u_mem/_0105_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold105 (.A(\u_ppwm/u_mem/memory[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold106 (.A(\u_ppwm/u_mem/_0071_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold107 (.A(\u_ppwm/u_mem/memory[88] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold108 (.A(\u_ppwm/u_mem/memory[61] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_ppwm/u_mem/memory[106] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold110 (.A(\u_ppwm/u_mem/_0112_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold111 (.A(\u_ppwm/u_mem/memory[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold112 (.A(\u_ppwm/u_mem/memory[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_ppwm/u_mem/_0050_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold114 (.A(\u_ppwm/u_mem/memory[98] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold115 (.A(\u_ppwm/u_mem/_0104_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold116 (.A(\u_ppwm/u_mem/memory[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold117 (.A(\u_ppwm/u_mem/memory[58] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold118 (.A(\u_ppwm/u_mem/_0064_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold119 (.A(\u_ppwm/u_mem/memory[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold120 (.A(\u_ppwm/u_mem/memory[102] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold121 (.A(\u_ppwm/u_mem/memory[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold122 (.A(\u_ppwm/u_mem/memory[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_ppwm/u_mem/_0044_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold124 (.A(\u_ppwm/u_mem/memory[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold125 (.A(\u_ppwm/u_mem/_0084_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold126 (.A(\u_ppwm/u_mem/memory[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_ppwm/u_mem/_0037_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_ppwm/u_mem/memory[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold129 (.A(\u_ppwm/u_mem/_0089_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_ppwm/u_mem/memory[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold131 (.A(\u_ppwm/u_mem/memory[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_ppwm/u_mem/_0035_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold133 (.A(\u_ppwm/u_mem/memory[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold134 (.A(\u_ppwm/u_mem/_0026_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold135 (.A(\u_ppwm/u_mem/state_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_ppwm/u_mem/_0004_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold137 (.A(\u_ppwm/u_mem/memory[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold138 (.A(\u_ppwm/u_mem/memory[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_ppwm/u_mem/memory[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold140 (.A(\u_ppwm/u_mem/_0043_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_ppwm/u_mem/memory[95] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold142 (.A(\u_ppwm/u_mem/_0101_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold143 (.A(\u_ppwm/u_mem/memory[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold144 (.A(\u_ppwm/u_mem/_0009_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_ppwm/u_mem/memory[105] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_ppwm/u_mem/_0111_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_ppwm/u_mem/memory[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold148 (.A(\u_ppwm/u_mem/_0082_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold149 (.A(\u_ppwm/u_mem/memory[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold150 (.A(\u_ppwm/u_mem/memory[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold151 (.A(\u_ppwm/u_mem/_0076_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_ppwm/u_mem/memory[94] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_ppwm/u_mem/_0100_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold154 (.A(\u_ppwm/u_mem/memory[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_ppwm/u_mem/_0049_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold156 (.A(\u_ppwm/u_mem/memory[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_ppwm/u_mem/_0029_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold158 (.A(\u_ppwm/u_mem/memory[92] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_ppwm/u_mem/_0001_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_ppwm/u_mem/memory[103] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold161 (.A(\u_ppwm/u_mem/memory[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_ppwm/u_mem/_0025_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold163 (.A(\u_ppwm/u_mem/memory[57] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold164 (.A(\u_ppwm/u_mem/memory[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold165 (.A(\u_ppwm/u_pwm/cmp_value[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold166 (.A(\u_ppwm/u_pwm/_003_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold167 (.A(\u_ppwm/u_mem/_0003_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold168 (.A(\u_ppwm/u_mem/memory[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_ppwm/u_mem/memory[104] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold170 (.A(\u_ppwm/u_mem/memory[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold171 (.A(\u_ppwm/u_mem/_0091_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold172 (.A(\u_ppwm/u_mem/memory[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold173 (.A(\u_ppwm/u_mem/memory[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold174 (.A(\u_ppwm/u_mem/memory[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold175 (.A(\u_ppwm/u_mem/memory[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_ppwm/u_mem/_0023_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold177 (.A(\u_ppwm/u_mem/memory[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold178 (.A(\u_ppwm/u_pwm/counter[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_ppwm/u_pwm/_028_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold180 (.A(\u_ppwm/u_pwm/_017_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_ppwm/u_pwm/counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold182 (.A(\u_ppwm/u_pwm/_011_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold183 (.A(\u_ppwm/u_mem/memory[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold184 (.A(\u_ppwm/u_mem/_0022_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold185 (.A(\u_ppwm/u_mem/memory[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_ppwm/u_mem/memory[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold187 (.A(\u_ppwm/u_mem/_0036_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold188 (.A(\u_ppwm/u_mem/memory[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_ppwm/u_mem/_0048_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold190 (.A(\u_ppwm/u_mem/memory[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold191 (.A(\u_ppwm/u_mem/memory[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold192 (.A(\u_ppwm/u_mem/memory[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_ppwm/u_mem/memory[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold194 (.A(\u_ppwm/u_mem/_0015_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_ppwm/u_mem/memory[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold196 (.A(\u_ppwm/u_mem/memory[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_ppwm/u_mem/bit_count[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold198 (.A(\u_ppwm/u_mem/_0489_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_ppwm/u_mem/_0125_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold200 (.A(\u_ppwm/u_mem/memory[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold201 (.A(\u_ppwm/u_mem/_0092_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold202 (.A(\u_ppwm/u_mem/memory[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold203 (.A(\u_ppwm/u_mem/memory[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold204 (.A(\u_ppwm/u_pwm/counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_ppwm/u_pwm/_101_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold206 (.A(\u_ppwm/u_pwm/_012_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold207 (.A(\u_ppwm/global_counter[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold208 (.A(\u_ppwm/u_global_counter/_010_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold209 (.A(\u_ppwm/u_mem/memory[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold210 (.A(\u_ppwm/u_mem/_0008_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold211 (.A(\u_ppwm/u_mem/memory[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold212 (.A(\u_ppwm/u_mem/memory[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold213 (.A(\u_ppwm/u_mem/memory[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold214 (.A(\u_ppwm/u_mem/memory[93] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold215 (.A(\u_ppwm/u_mem/memory[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold216 (.A(\u_ppwm/u_mem/_0083_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold217 (.A(\u_ppwm/global_counter[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold218 (.A(\u_ppwm/u_global_counter/_019_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold219 (.A(\u_ppwm/u_mem/bit_count[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold220 (.A(\u_ppwm/u_mem/_0487_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold221 (.A(\u_ppwm/u_mem/_0124_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold222 (.A(\u_ppwm/global_counter[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_ppwm/u_global_counter/_004_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold224 (.A(\u_ppwm/u_mem/memory[62] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold225 (.A(\u_ppwm/u_pwm/counter[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold226 (.A(\u_ppwm/u_pwm/_033_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold227 (.A(\u_ppwm/u_pwm/_020_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold228 (.A(\u_ppwm/u_mem/memory[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold229 (.A(\u_ppwm/u_mem/memory[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold230 (.A(\u_ppwm/u_mem/_0007_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold231 (.A(\u_ppwm/global_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_ppwm/u_global_counter/_003_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold233 (.A(\u_ppwm/u_pwm/counter[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold234 (.A(\u_ppwm/u_pwm/_025_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold235 (.A(\u_ppwm/u_pwm/_015_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold236 (.A(\u_ppwm/global_counter[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold237 (.A(\u_ppwm/u_global_counter/_006_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold238 (.A(\u_ppwm/u_mem/bit_count[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold239 (.A(\u_ppwm/u_mem/_0483_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold240 (.A(\u_ppwm/global_counter[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold241 (.A(\u_ppwm/u_global_counter/_045_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold242 (.A(\u_ppwm/u_global_counter/_014_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold243 (.A(\u_ppwm/u_mem/bit_count[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold244 (.A(\u_ppwm/u_mem/_0481_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold245 (.A(\u_ppwm/u_mem/_0121_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold246 (.A(\u_ppwm/u_ex/state_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold247 (.A(\u_ppwm/u_ex/_0055_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold248 (.A(\u_ppwm/u_ex/_0000_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold249 (.A(\u_ppwm/u_mem/bit_count[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold250 (.A(\u_ppwm/u_mem/bit_count[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold251 (.A(\u_ppwm/u_mem/_0247_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold252 (.A(\u_ppwm/global_counter[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold253 (.A(\u_ppwm/u_global_counter/_018_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold254 (.A(\u_ppwm/global_counter[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold255 (.A(\u_ppwm/u_global_counter/_015_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold256 (.A(\u_ppwm/u_mem/bit_count[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold257 (.A(\u_ppwm/mem_write_done ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold258 (.A(\u_ppwm/u_mem/_0005_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold259 (.A(\u_ppwm/global_counter[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold260 (.A(\u_ppwm/u_global_counter/_033_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold261 (.A(\u_ppwm/u_global_counter/_005_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold262 (.A(\u_ppwm/global_counter[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold263 (.A(\u_ppwm/u_global_counter/_036_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold264 (.A(\u_ppwm/u_global_counter/_007_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold265 (.A(\u_ppwm/global_counter[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold266 (.A(\u_ppwm/u_global_counter/_043_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold267 (.A(\u_ppwm/u_global_counter/_013_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold268 (.A(\u_ppwm/u_pwm/counter[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold269 (.A(\u_ppwm/u_pwm/_029_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold270 (.A(\u_ppwm/u_mem/bit_count[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold271 (.A(\u_ppwm/global_counter[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold272 (.A(\u_ppwm/u_global_counter/_039_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold273 (.A(\u_ppwm/u_global_counter/_011_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold274 (.A(\u_ppwm/period_start ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold275 (.A(\u_ppwm/u_ex/_0002_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold276 (.A(\u_ppwm/u_pwm/counter[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold277 (.A(\u_ppwm/global_counter[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold278 (.A(\u_ppwm/u_global_counter/_017_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold279 (.A(\u_ppwm/u_pwm/counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold280 (.A(\u_ppwm/u_ex/cmp_flag_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold281 (.A(\u_ppwm/u_ex/_0216_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold282 (.A(\u_ppwm/u_ex/_0007_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold283 (.A(\u_ppwm/u_pwm/counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold284 (.A(\u_ppwm/u_pwm/counter[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold285 (.A(\u_ppwm/global_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold286 (.A(\u_ppwm/global_counter[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold287 (.A(\u_ppwm/global_counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold288 (.A(\u_ppwm/u_global_counter/_002_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold289 (.A(\u_ppwm/u_ex/reg_value_q[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold290 (.A(\u_ppwm/u_ex/_0028_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold291 (.A(\u_ppwm/global_counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold292 (.A(\u_ppwm/u_ex/reg_value_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold293 (.A(\u_ppwm/u_ex/_0009_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold294 (.A(\u_ppwm/u_ex/reg_value_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_ppwm/u_ex/reg_value_q[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold296 (.A(\u_ppwm/pwm_value[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold297 (.A(\u_ppwm/global_counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold298 (.A(\u_ppwm/u_global_counter/_034_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold299 (.A(\u_ppwm/u_ex/reg_value_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold300 (.A(\u_ppwm/u_ex/reg_value_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold301 (.A(\u_ppwm/pwm_value[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold302 (.A(\u_ppwm/u_ex/_0014_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold303 (.A(\u_ppwm/u_ex/reg_value_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold304 (.A(\u_ppwm/pwm_value[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold305 (.A(\u_ppwm/pc[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold306 (.A(\u_ppwm/u_ex/_0078_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold307 (.A(\u_ppwm/pwm_value[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold308 (.A(\u_ppwm/pwm_value[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold309 (.A(\u_ppwm/pwm_value[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold310 (.A(\u_ppwm/u_ex/reg_value_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold311 (.A(\u_ppwm/u_ex/_0020_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold312 (.A(\u_ppwm/pwm_value[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold313 (.A(\u_ppwm/u_ex/reg_value_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold314 (.A(\u_ppwm/u_ex/reg_value_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold315 (.A(\u_ppwm/pc[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold316 (.A(\u_ppwm/u_ex/_0086_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold317 (.A(\u_ppwm/u_ex/_0006_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold318 (.A(\u_ppwm/u_ex/state_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold319 (.A(\u_ppwm/pwm_value[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold320 (.A(\u_ppwm/u_ex/_0010_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold321 (.A(\u_ppwm/pc[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold322 (.A(\u_ppwm/pwm_value[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold323 (.A(\u_ppwm/u_mem/bit_count[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold324 (.A(\u_ppwm/pwm_value[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net692));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
 assign uo_out[1] = net19;
 assign uo_out[2] = net20;
 assign uo_out[3] = net21;
 assign uo_out[4] = net22;
 assign uo_out[5] = net23;
 assign uo_out[6] = net24;
 assign uo_out[7] = net25;
endmodule
