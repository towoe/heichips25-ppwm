module heichips25_ppwm (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire \u_ppwm/global_counter_high[0] ;
 wire \u_ppwm/global_counter_high[10] ;
 wire \u_ppwm/global_counter_high[11] ;
 wire \u_ppwm/global_counter_high[12] ;
 wire \u_ppwm/global_counter_high[13] ;
 wire \u_ppwm/global_counter_high[14] ;
 wire \u_ppwm/global_counter_high[15] ;
 wire \u_ppwm/global_counter_high[16] ;
 wire \u_ppwm/global_counter_high[17] ;
 wire \u_ppwm/global_counter_high[18] ;
 wire \u_ppwm/global_counter_high[19] ;
 wire \u_ppwm/global_counter_high[1] ;
 wire \u_ppwm/global_counter_high[2] ;
 wire \u_ppwm/global_counter_high[3] ;
 wire \u_ppwm/global_counter_high[4] ;
 wire \u_ppwm/global_counter_high[5] ;
 wire \u_ppwm/global_counter_high[6] ;
 wire \u_ppwm/global_counter_high[7] ;
 wire \u_ppwm/global_counter_high[8] ;
 wire \u_ppwm/global_counter_high[9] ;
 wire \u_ppwm/instr[0] ;
 wire \u_ppwm/instr[1] ;
 wire \u_ppwm/instr[2] ;
 wire \u_ppwm/instr[3] ;
 wire \u_ppwm/instr[4] ;
 wire \u_ppwm/instr[5] ;
 wire \u_ppwm/instr[6] ;
 wire \u_ppwm/mem_write_done ;
 wire \u_ppwm/pc[0] ;
 wire \u_ppwm/pc[1] ;
 wire \u_ppwm/pc[2] ;
 wire \u_ppwm/pc[3] ;
 wire \u_ppwm/period_start ;
 wire \u_ppwm/pwm_value[0] ;
 wire \u_ppwm/pwm_value[1] ;
 wire \u_ppwm/pwm_value[2] ;
 wire \u_ppwm/pwm_value[3] ;
 wire \u_ppwm/pwm_value[4] ;
 wire \u_ppwm/pwm_value[5] ;
 wire \u_ppwm/pwm_value[6] ;
 wire \u_ppwm/pwm_value[7] ;
 wire \u_ppwm/pwm_value[8] ;
 wire \u_ppwm/pwm_value[9] ;
 wire \u_ppwm/u_ex/_000_ ;
 wire \u_ppwm/u_ex/_001_ ;
 wire \u_ppwm/u_ex/_002_ ;
 wire \u_ppwm/u_ex/_003_ ;
 wire \u_ppwm/u_ex/_004_ ;
 wire \u_ppwm/u_ex/_005_ ;
 wire \u_ppwm/u_ex/_006_ ;
 wire \u_ppwm/u_ex/_007_ ;
 wire \u_ppwm/u_ex/_008_ ;
 wire \u_ppwm/u_ex/_009_ ;
 wire \u_ppwm/u_ex/_010_ ;
 wire \u_ppwm/u_ex/_011_ ;
 wire \u_ppwm/u_ex/_012_ ;
 wire \u_ppwm/u_ex/_013_ ;
 wire \u_ppwm/u_ex/_014_ ;
 wire \u_ppwm/u_ex/_015_ ;
 wire \u_ppwm/u_ex/_016_ ;
 wire \u_ppwm/u_ex/_017_ ;
 wire \u_ppwm/u_ex/_018_ ;
 wire \u_ppwm/u_ex/_019_ ;
 wire \u_ppwm/u_ex/_020_ ;
 wire \u_ppwm/u_ex/_021_ ;
 wire \u_ppwm/u_ex/_022_ ;
 wire \u_ppwm/u_ex/_023_ ;
 wire \u_ppwm/u_ex/_024_ ;
 wire \u_ppwm/u_ex/_025_ ;
 wire \u_ppwm/u_ex/_026_ ;
 wire \u_ppwm/u_ex/_027_ ;
 wire \u_ppwm/u_ex/_028_ ;
 wire \u_ppwm/u_ex/_029_ ;
 wire \u_ppwm/u_ex/_030_ ;
 wire \u_ppwm/u_ex/_031_ ;
 wire \u_ppwm/u_ex/_032_ ;
 wire \u_ppwm/u_ex/_033_ ;
 wire \u_ppwm/u_ex/_034_ ;
 wire \u_ppwm/u_ex/_035_ ;
 wire \u_ppwm/u_ex/_036_ ;
 wire \u_ppwm/u_ex/_037_ ;
 wire \u_ppwm/u_ex/_038_ ;
 wire \u_ppwm/u_ex/_039_ ;
 wire \u_ppwm/u_ex/_040_ ;
 wire \u_ppwm/u_ex/_041_ ;
 wire \u_ppwm/u_ex/_042_ ;
 wire \u_ppwm/u_ex/_043_ ;
 wire \u_ppwm/u_ex/_044_ ;
 wire \u_ppwm/u_ex/_045_ ;
 wire \u_ppwm/u_ex/_046_ ;
 wire \u_ppwm/u_ex/_047_ ;
 wire \u_ppwm/u_ex/_048_ ;
 wire \u_ppwm/u_ex/_049_ ;
 wire \u_ppwm/u_ex/_050_ ;
 wire \u_ppwm/u_ex/_051_ ;
 wire \u_ppwm/u_ex/_052_ ;
 wire \u_ppwm/u_ex/_053_ ;
 wire \u_ppwm/u_ex/_054_ ;
 wire \u_ppwm/u_ex/_055_ ;
 wire \u_ppwm/u_ex/_056_ ;
 wire \u_ppwm/u_ex/_057_ ;
 wire \u_ppwm/u_ex/_058_ ;
 wire \u_ppwm/u_ex/_059_ ;
 wire \u_ppwm/u_ex/_060_ ;
 wire \u_ppwm/u_ex/_061_ ;
 wire \u_ppwm/u_ex/_062_ ;
 wire \u_ppwm/u_ex/_063_ ;
 wire \u_ppwm/u_ex/_064_ ;
 wire \u_ppwm/u_ex/_065_ ;
 wire \u_ppwm/u_ex/_066_ ;
 wire \u_ppwm/u_ex/_067_ ;
 wire \u_ppwm/u_ex/_068_ ;
 wire \u_ppwm/u_ex/_069_ ;
 wire \u_ppwm/u_ex/_070_ ;
 wire \u_ppwm/u_ex/_071_ ;
 wire \u_ppwm/u_ex/_072_ ;
 wire \u_ppwm/u_ex/_073_ ;
 wire \u_ppwm/u_ex/_074_ ;
 wire \u_ppwm/u_ex/_075_ ;
 wire \u_ppwm/u_ex/_076_ ;
 wire \u_ppwm/u_ex/_077_ ;
 wire \u_ppwm/u_ex/_078_ ;
 wire \u_ppwm/u_ex/_079_ ;
 wire \u_ppwm/u_ex/_080_ ;
 wire \u_ppwm/u_ex/_081_ ;
 wire \u_ppwm/u_ex/_082_ ;
 wire \u_ppwm/u_ex/_083_ ;
 wire \u_ppwm/u_ex/_084_ ;
 wire \u_ppwm/u_ex/_085_ ;
 wire \u_ppwm/u_ex/_086_ ;
 wire \u_ppwm/u_ex/_087_ ;
 wire \u_ppwm/u_ex/_088_ ;
 wire \u_ppwm/u_ex/_089_ ;
 wire \u_ppwm/u_ex/_090_ ;
 wire \u_ppwm/u_ex/_091_ ;
 wire \u_ppwm/u_ex/_092_ ;
 wire \u_ppwm/u_ex/_093_ ;
 wire \u_ppwm/u_ex/_094_ ;
 wire \u_ppwm/u_ex/_095_ ;
 wire \u_ppwm/u_ex/_096_ ;
 wire \u_ppwm/u_ex/_097_ ;
 wire \u_ppwm/u_ex/_098_ ;
 wire \u_ppwm/u_ex/_099_ ;
 wire \u_ppwm/u_ex/_100_ ;
 wire \u_ppwm/u_ex/_101_ ;
 wire \u_ppwm/u_ex/_102_ ;
 wire \u_ppwm/u_ex/_103_ ;
 wire \u_ppwm/u_ex/_104_ ;
 wire \u_ppwm/u_ex/_105_ ;
 wire \u_ppwm/u_ex/_106_ ;
 wire \u_ppwm/u_ex/_107_ ;
 wire \u_ppwm/u_ex/_108_ ;
 wire \u_ppwm/u_ex/_109_ ;
 wire \u_ppwm/u_ex/_110_ ;
 wire \u_ppwm/u_ex/_111_ ;
 wire \u_ppwm/u_ex/_112_ ;
 wire \u_ppwm/u_ex/_113_ ;
 wire \u_ppwm/u_ex/_114_ ;
 wire \u_ppwm/u_ex/_115_ ;
 wire \u_ppwm/u_ex/_116_ ;
 wire \u_ppwm/u_ex/_117_ ;
 wire \u_ppwm/u_ex/_118_ ;
 wire \u_ppwm/u_ex/_119_ ;
 wire \u_ppwm/u_ex/_120_ ;
 wire \u_ppwm/u_ex/_121_ ;
 wire \u_ppwm/u_ex/_122_ ;
 wire \u_ppwm/u_ex/_123_ ;
 wire \u_ppwm/u_ex/_124_ ;
 wire \u_ppwm/u_ex/_125_ ;
 wire \u_ppwm/u_ex/_126_ ;
 wire \u_ppwm/u_ex/_127_ ;
 wire \u_ppwm/u_ex/_128_ ;
 wire \u_ppwm/u_ex/_129_ ;
 wire \u_ppwm/u_ex/_130_ ;
 wire \u_ppwm/u_ex/_131_ ;
 wire \u_ppwm/u_ex/_132_ ;
 wire \u_ppwm/u_ex/_133_ ;
 wire \u_ppwm/u_ex/_134_ ;
 wire \u_ppwm/u_ex/_135_ ;
 wire \u_ppwm/u_ex/_136_ ;
 wire \u_ppwm/u_ex/_137_ ;
 wire \u_ppwm/u_ex/_138_ ;
 wire \u_ppwm/u_ex/_139_ ;
 wire \u_ppwm/u_ex/_140_ ;
 wire \u_ppwm/u_ex/_141_ ;
 wire \u_ppwm/u_ex/_142_ ;
 wire \u_ppwm/u_ex/_143_ ;
 wire \u_ppwm/u_ex/_144_ ;
 wire \u_ppwm/u_ex/_145_ ;
 wire \u_ppwm/u_ex/_146_ ;
 wire \u_ppwm/u_ex/_147_ ;
 wire \u_ppwm/u_ex/_148_ ;
 wire \u_ppwm/u_ex/_149_ ;
 wire \u_ppwm/u_ex/_150_ ;
 wire \u_ppwm/u_ex/_151_ ;
 wire \u_ppwm/u_ex/_152_ ;
 wire \u_ppwm/u_ex/_153_ ;
 wire \u_ppwm/u_ex/_154_ ;
 wire \u_ppwm/u_ex/_155_ ;
 wire \u_ppwm/u_ex/_156_ ;
 wire \u_ppwm/u_ex/_157_ ;
 wire \u_ppwm/u_ex/_158_ ;
 wire \u_ppwm/u_ex/_159_ ;
 wire \u_ppwm/u_ex/_160_ ;
 wire \u_ppwm/u_ex/_161_ ;
 wire \u_ppwm/u_ex/_162_ ;
 wire \u_ppwm/u_ex/_163_ ;
 wire \u_ppwm/u_ex/_164_ ;
 wire \u_ppwm/u_ex/_165_ ;
 wire \u_ppwm/u_ex/_166_ ;
 wire \u_ppwm/u_ex/_167_ ;
 wire \u_ppwm/u_ex/_168_ ;
 wire \u_ppwm/u_ex/_169_ ;
 wire \u_ppwm/u_ex/_170_ ;
 wire \u_ppwm/u_ex/_171_ ;
 wire \u_ppwm/u_ex/_172_ ;
 wire \u_ppwm/u_ex/_173_ ;
 wire \u_ppwm/u_ex/_174_ ;
 wire \u_ppwm/u_ex/_175_ ;
 wire \u_ppwm/u_ex/_176_ ;
 wire \u_ppwm/u_ex/_177_ ;
 wire \u_ppwm/u_ex/_178_ ;
 wire \u_ppwm/u_ex/_179_ ;
 wire \u_ppwm/u_ex/_180_ ;
 wire \u_ppwm/u_ex/_181_ ;
 wire \u_ppwm/u_ex/_182_ ;
 wire \u_ppwm/u_ex/_183_ ;
 wire \u_ppwm/u_ex/_184_ ;
 wire \u_ppwm/u_ex/_185_ ;
 wire \u_ppwm/u_ex/_186_ ;
 wire \u_ppwm/u_ex/_187_ ;
 wire \u_ppwm/u_ex/_188_ ;
 wire \u_ppwm/u_ex/_189_ ;
 wire \u_ppwm/u_ex/_190_ ;
 wire \u_ppwm/u_ex/_191_ ;
 wire \u_ppwm/u_ex/_192_ ;
 wire \u_ppwm/u_ex/_193_ ;
 wire \u_ppwm/u_ex/_194_ ;
 wire \u_ppwm/u_ex/_195_ ;
 wire \u_ppwm/u_ex/_196_ ;
 wire \u_ppwm/u_ex/_197_ ;
 wire \u_ppwm/u_ex/_198_ ;
 wire \u_ppwm/u_ex/_199_ ;
 wire \u_ppwm/u_ex/_200_ ;
 wire \u_ppwm/u_ex/_201_ ;
 wire \u_ppwm/u_ex/_202_ ;
 wire \u_ppwm/u_ex/_203_ ;
 wire \u_ppwm/u_ex/_204_ ;
 wire \u_ppwm/u_ex/_205_ ;
 wire \u_ppwm/u_ex/_206_ ;
 wire \u_ppwm/u_ex/_207_ ;
 wire \u_ppwm/u_ex/_208_ ;
 wire \u_ppwm/u_ex/_209_ ;
 wire \u_ppwm/u_ex/_210_ ;
 wire \u_ppwm/u_ex/_211_ ;
 wire \u_ppwm/u_ex/_212_ ;
 wire \u_ppwm/u_ex/_213_ ;
 wire \u_ppwm/u_ex/_214_ ;
 wire \u_ppwm/u_ex/_215_ ;
 wire \u_ppwm/u_ex/_216_ ;
 wire \u_ppwm/u_ex/_217_ ;
 wire \u_ppwm/u_ex/_218_ ;
 wire \u_ppwm/u_ex/_219_ ;
 wire \u_ppwm/u_ex/_220_ ;
 wire \u_ppwm/u_ex/_221_ ;
 wire \u_ppwm/u_ex/_222_ ;
 wire \u_ppwm/u_ex/_223_ ;
 wire \u_ppwm/u_ex/_224_ ;
 wire \u_ppwm/u_ex/_225_ ;
 wire \u_ppwm/u_ex/_226_ ;
 wire \u_ppwm/u_ex/_227_ ;
 wire \u_ppwm/u_ex/_228_ ;
 wire \u_ppwm/u_ex/_229_ ;
 wire \u_ppwm/u_ex/_230_ ;
 wire \u_ppwm/u_ex/_231_ ;
 wire \u_ppwm/u_ex/_232_ ;
 wire \u_ppwm/u_ex/_233_ ;
 wire \u_ppwm/u_ex/_234_ ;
 wire \u_ppwm/u_ex/_235_ ;
 wire \u_ppwm/u_ex/_236_ ;
 wire \u_ppwm/u_ex/_237_ ;
 wire \u_ppwm/u_ex/_238_ ;
 wire \u_ppwm/u_ex/_239_ ;
 wire \u_ppwm/u_ex/_240_ ;
 wire \u_ppwm/u_ex/_241_ ;
 wire \u_ppwm/u_ex/_242_ ;
 wire \u_ppwm/u_ex/_243_ ;
 wire \u_ppwm/u_ex/_244_ ;
 wire \u_ppwm/u_ex/_245_ ;
 wire \u_ppwm/u_ex/_246_ ;
 wire \u_ppwm/u_ex/_247_ ;
 wire \u_ppwm/u_ex/_248_ ;
 wire \u_ppwm/u_ex/_249_ ;
 wire \u_ppwm/u_ex/_250_ ;
 wire \u_ppwm/u_ex/_251_ ;
 wire \u_ppwm/u_ex/_252_ ;
 wire \u_ppwm/u_ex/_253_ ;
 wire \u_ppwm/u_ex/_254_ ;
 wire \u_ppwm/u_ex/_255_ ;
 wire \u_ppwm/u_ex/_256_ ;
 wire \u_ppwm/u_ex/_257_ ;
 wire \u_ppwm/u_ex/_258_ ;
 wire \u_ppwm/u_ex/_259_ ;
 wire \u_ppwm/u_ex/_260_ ;
 wire \u_ppwm/u_ex/_261_ ;
 wire \u_ppwm/u_ex/_262_ ;
 wire \u_ppwm/u_ex/_263_ ;
 wire \u_ppwm/u_ex/_264_ ;
 wire \u_ppwm/u_ex/_265_ ;
 wire \u_ppwm/u_ex/_266_ ;
 wire \u_ppwm/u_ex/_267_ ;
 wire \u_ppwm/u_ex/_268_ ;
 wire \u_ppwm/u_ex/_269_ ;
 wire \u_ppwm/u_ex/_270_ ;
 wire \u_ppwm/u_ex/_271_ ;
 wire \u_ppwm/u_ex/_272_ ;
 wire \u_ppwm/u_ex/_273_ ;
 wire \u_ppwm/u_ex/_274_ ;
 wire \u_ppwm/u_ex/_275_ ;
 wire \u_ppwm/u_ex/_276_ ;
 wire \u_ppwm/u_ex/_277_ ;
 wire \u_ppwm/u_ex/_278_ ;
 wire \u_ppwm/u_ex/_279_ ;
 wire \u_ppwm/u_ex/_280_ ;
 wire \u_ppwm/u_ex/_281_ ;
 wire \u_ppwm/u_ex/_282_ ;
 wire \u_ppwm/u_ex/_283_ ;
 wire \u_ppwm/u_ex/_284_ ;
 wire \u_ppwm/u_ex/_285_ ;
 wire \u_ppwm/u_ex/_286_ ;
 wire \u_ppwm/u_ex/_287_ ;
 wire \u_ppwm/u_ex/_288_ ;
 wire \u_ppwm/u_ex/_289_ ;
 wire \u_ppwm/u_ex/_290_ ;
 wire \u_ppwm/u_ex/_291_ ;
 wire \u_ppwm/u_ex/_292_ ;
 wire \u_ppwm/u_ex/_293_ ;
 wire \u_ppwm/u_ex/_294_ ;
 wire \u_ppwm/u_ex/_295_ ;
 wire \u_ppwm/u_ex/_296_ ;
 wire \u_ppwm/u_ex/_297_ ;
 wire \u_ppwm/u_ex/_298_ ;
 wire \u_ppwm/u_ex/_299_ ;
 wire \u_ppwm/u_ex/_300_ ;
 wire \u_ppwm/u_ex/_301_ ;
 wire \u_ppwm/u_ex/_302_ ;
 wire \u_ppwm/u_ex/_303_ ;
 wire \u_ppwm/u_ex/_304_ ;
 wire \u_ppwm/u_ex/_305_ ;
 wire \u_ppwm/u_ex/_306_ ;
 wire \u_ppwm/u_ex/_307_ ;
 wire \u_ppwm/u_ex/_308_ ;
 wire \u_ppwm/u_ex/_309_ ;
 wire \u_ppwm/u_ex/_310_ ;
 wire \u_ppwm/u_ex/_311_ ;
 wire \u_ppwm/u_ex/_312_ ;
 wire \u_ppwm/u_ex/_313_ ;
 wire \u_ppwm/u_ex/_314_ ;
 wire \u_ppwm/u_ex/_315_ ;
 wire \u_ppwm/u_ex/_316_ ;
 wire \u_ppwm/u_ex/_317_ ;
 wire \u_ppwm/u_ex/_318_ ;
 wire \u_ppwm/u_ex/_319_ ;
 wire \u_ppwm/u_ex/_320_ ;
 wire \u_ppwm/u_ex/_321_ ;
 wire \u_ppwm/u_ex/_322_ ;
 wire \u_ppwm/u_ex/_323_ ;
 wire \u_ppwm/u_ex/_324_ ;
 wire \u_ppwm/u_ex/_325_ ;
 wire \u_ppwm/u_ex/_326_ ;
 wire \u_ppwm/u_ex/_327_ ;
 wire \u_ppwm/u_ex/_328_ ;
 wire \u_ppwm/u_ex/_329_ ;
 wire \u_ppwm/u_ex/_330_ ;
 wire \u_ppwm/u_ex/_331_ ;
 wire \u_ppwm/u_ex/_332_ ;
 wire \u_ppwm/u_ex/_333_ ;
 wire \u_ppwm/u_ex/_334_ ;
 wire \u_ppwm/u_ex/_335_ ;
 wire \u_ppwm/u_ex/_336_ ;
 wire \u_ppwm/u_ex/_337_ ;
 wire \u_ppwm/u_ex/_338_ ;
 wire \u_ppwm/u_ex/_339_ ;
 wire \u_ppwm/u_ex/_340_ ;
 wire \u_ppwm/u_ex/_341_ ;
 wire \u_ppwm/u_ex/_342_ ;
 wire \u_ppwm/u_ex/_343_ ;
 wire \u_ppwm/u_ex/_344_ ;
 wire \u_ppwm/u_ex/_345_ ;
 wire \u_ppwm/u_ex/_346_ ;
 wire \u_ppwm/u_ex/_347_ ;
 wire \u_ppwm/u_ex/_348_ ;
 wire \u_ppwm/u_ex/_349_ ;
 wire \u_ppwm/u_ex/_350_ ;
 wire \u_ppwm/u_ex/_351_ ;
 wire \u_ppwm/u_ex/_352_ ;
 wire \u_ppwm/u_ex/_353_ ;
 wire \u_ppwm/u_ex/_354_ ;
 wire \u_ppwm/u_ex/_355_ ;
 wire \u_ppwm/u_ex/_356_ ;
 wire \u_ppwm/u_ex/_357_ ;
 wire \u_ppwm/u_ex/_358_ ;
 wire \u_ppwm/u_ex/_359_ ;
 wire \u_ppwm/u_ex/_360_ ;
 wire \u_ppwm/u_ex/_361_ ;
 wire \u_ppwm/u_ex/_362_ ;
 wire \u_ppwm/u_ex/_363_ ;
 wire \u_ppwm/u_ex/_364_ ;
 wire \u_ppwm/u_ex/_365_ ;
 wire \u_ppwm/u_ex/_366_ ;
 wire \u_ppwm/u_ex/_367_ ;
 wire \u_ppwm/u_ex/_368_ ;
 wire \u_ppwm/u_ex/_369_ ;
 wire \u_ppwm/u_ex/_370_ ;
 wire \u_ppwm/u_ex/_371_ ;
 wire \u_ppwm/u_ex/_372_ ;
 wire \u_ppwm/u_ex/_373_ ;
 wire \u_ppwm/u_ex/_374_ ;
 wire \u_ppwm/u_ex/_375_ ;
 wire \u_ppwm/u_ex/_376_ ;
 wire \u_ppwm/u_ex/_377_ ;
 wire \u_ppwm/u_ex/_378_ ;
 wire \u_ppwm/u_ex/_379_ ;
 wire \u_ppwm/u_ex/_380_ ;
 wire \u_ppwm/u_ex/_381_ ;
 wire \u_ppwm/u_ex/_382_ ;
 wire \u_ppwm/u_ex/_383_ ;
 wire \u_ppwm/u_ex/_384_ ;
 wire \u_ppwm/u_ex/_385_ ;
 wire \u_ppwm/u_ex/_386_ ;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire \u_ppwm/u_ex/cmp_flag_q ;
 wire \u_ppwm/u_ex/reg_value_q[0] ;
 wire \u_ppwm/u_ex/reg_value_q[1] ;
 wire \u_ppwm/u_ex/reg_value_q[2] ;
 wire \u_ppwm/u_ex/reg_value_q[3] ;
 wire \u_ppwm/u_ex/reg_value_q[4] ;
 wire \u_ppwm/u_ex/reg_value_q[5] ;
 wire \u_ppwm/u_ex/reg_value_q[6] ;
 wire \u_ppwm/u_ex/reg_value_q[7] ;
 wire \u_ppwm/u_ex/reg_value_q[8] ;
 wire \u_ppwm/u_ex/reg_value_q[9] ;
 wire \u_ppwm/u_ex/state_q[0] ;
 wire \u_ppwm/u_ex/state_q[1] ;
 wire \u_ppwm/u_ex/state_q[2] ;
 wire \u_ppwm/u_global_counter/_000_ ;
 wire \u_ppwm/u_global_counter/_001_ ;
 wire \u_ppwm/u_global_counter/_002_ ;
 wire \u_ppwm/u_global_counter/_003_ ;
 wire \u_ppwm/u_global_counter/_004_ ;
 wire \u_ppwm/u_global_counter/_005_ ;
 wire \u_ppwm/u_global_counter/_006_ ;
 wire \u_ppwm/u_global_counter/_007_ ;
 wire \u_ppwm/u_global_counter/_008_ ;
 wire \u_ppwm/u_global_counter/_009_ ;
 wire \u_ppwm/u_global_counter/_010_ ;
 wire \u_ppwm/u_global_counter/_011_ ;
 wire \u_ppwm/u_global_counter/_012_ ;
 wire \u_ppwm/u_global_counter/_013_ ;
 wire \u_ppwm/u_global_counter/_014_ ;
 wire \u_ppwm/u_global_counter/_015_ ;
 wire \u_ppwm/u_global_counter/_016_ ;
 wire \u_ppwm/u_global_counter/_017_ ;
 wire \u_ppwm/u_global_counter/_018_ ;
 wire \u_ppwm/u_global_counter/_019_ ;
 wire \u_ppwm/u_global_counter/_020_ ;
 wire \u_ppwm/u_global_counter/_021_ ;
 wire \u_ppwm/u_global_counter/_022_ ;
 wire \u_ppwm/u_global_counter/_023_ ;
 wire \u_ppwm/u_global_counter/_024_ ;
 wire \u_ppwm/u_global_counter/_025_ ;
 wire \u_ppwm/u_global_counter/_026_ ;
 wire \u_ppwm/u_global_counter/_027_ ;
 wire \u_ppwm/u_global_counter/_028_ ;
 wire \u_ppwm/u_global_counter/_029_ ;
 wire \u_ppwm/u_global_counter/_030_ ;
 wire \u_ppwm/u_global_counter/_031_ ;
 wire \u_ppwm/u_global_counter/_032_ ;
 wire \u_ppwm/u_global_counter/_033_ ;
 wire \u_ppwm/u_global_counter/_034_ ;
 wire \u_ppwm/u_global_counter/_035_ ;
 wire \u_ppwm/u_global_counter/_036_ ;
 wire \u_ppwm/u_global_counter/_037_ ;
 wire \u_ppwm/u_global_counter/_038_ ;
 wire \u_ppwm/u_global_counter/_039_ ;
 wire \u_ppwm/u_global_counter/_040_ ;
 wire \u_ppwm/u_global_counter/_041_ ;
 wire \u_ppwm/u_global_counter/_042_ ;
 wire \u_ppwm/u_global_counter/_043_ ;
 wire \u_ppwm/u_global_counter/_044_ ;
 wire \u_ppwm/u_global_counter/_045_ ;
 wire \u_ppwm/u_global_counter/_046_ ;
 wire \u_ppwm/u_global_counter/_047_ ;
 wire \u_ppwm/u_global_counter/_048_ ;
 wire \u_ppwm/u_global_counter/_049_ ;
 wire \u_ppwm/u_global_counter/_050_ ;
 wire \u_ppwm/u_global_counter/_051_ ;
 wire \u_ppwm/u_global_counter/_052_ ;
 wire \u_ppwm/u_mem/_0000_ ;
 wire \u_ppwm/u_mem/_0001_ ;
 wire \u_ppwm/u_mem/_0002_ ;
 wire \u_ppwm/u_mem/_0003_ ;
 wire \u_ppwm/u_mem/_0004_ ;
 wire \u_ppwm/u_mem/_0005_ ;
 wire \u_ppwm/u_mem/_0006_ ;
 wire \u_ppwm/u_mem/_0007_ ;
 wire \u_ppwm/u_mem/_0008_ ;
 wire \u_ppwm/u_mem/_0009_ ;
 wire \u_ppwm/u_mem/_0010_ ;
 wire \u_ppwm/u_mem/_0011_ ;
 wire \u_ppwm/u_mem/_0012_ ;
 wire \u_ppwm/u_mem/_0013_ ;
 wire \u_ppwm/u_mem/_0014_ ;
 wire \u_ppwm/u_mem/_0015_ ;
 wire \u_ppwm/u_mem/_0016_ ;
 wire \u_ppwm/u_mem/_0017_ ;
 wire \u_ppwm/u_mem/_0018_ ;
 wire \u_ppwm/u_mem/_0019_ ;
 wire \u_ppwm/u_mem/_0020_ ;
 wire \u_ppwm/u_mem/_0021_ ;
 wire \u_ppwm/u_mem/_0022_ ;
 wire \u_ppwm/u_mem/_0023_ ;
 wire \u_ppwm/u_mem/_0024_ ;
 wire \u_ppwm/u_mem/_0025_ ;
 wire \u_ppwm/u_mem/_0026_ ;
 wire \u_ppwm/u_mem/_0027_ ;
 wire \u_ppwm/u_mem/_0028_ ;
 wire \u_ppwm/u_mem/_0029_ ;
 wire \u_ppwm/u_mem/_0030_ ;
 wire \u_ppwm/u_mem/_0031_ ;
 wire \u_ppwm/u_mem/_0032_ ;
 wire \u_ppwm/u_mem/_0033_ ;
 wire \u_ppwm/u_mem/_0034_ ;
 wire \u_ppwm/u_mem/_0035_ ;
 wire \u_ppwm/u_mem/_0036_ ;
 wire \u_ppwm/u_mem/_0037_ ;
 wire \u_ppwm/u_mem/_0038_ ;
 wire \u_ppwm/u_mem/_0039_ ;
 wire \u_ppwm/u_mem/_0040_ ;
 wire \u_ppwm/u_mem/_0041_ ;
 wire \u_ppwm/u_mem/_0042_ ;
 wire \u_ppwm/u_mem/_0043_ ;
 wire \u_ppwm/u_mem/_0044_ ;
 wire \u_ppwm/u_mem/_0045_ ;
 wire \u_ppwm/u_mem/_0046_ ;
 wire \u_ppwm/u_mem/_0047_ ;
 wire \u_ppwm/u_mem/_0048_ ;
 wire \u_ppwm/u_mem/_0049_ ;
 wire \u_ppwm/u_mem/_0050_ ;
 wire \u_ppwm/u_mem/_0051_ ;
 wire \u_ppwm/u_mem/_0052_ ;
 wire \u_ppwm/u_mem/_0053_ ;
 wire \u_ppwm/u_mem/_0054_ ;
 wire \u_ppwm/u_mem/_0055_ ;
 wire \u_ppwm/u_mem/_0056_ ;
 wire \u_ppwm/u_mem/_0057_ ;
 wire \u_ppwm/u_mem/_0058_ ;
 wire \u_ppwm/u_mem/_0059_ ;
 wire \u_ppwm/u_mem/_0060_ ;
 wire \u_ppwm/u_mem/_0061_ ;
 wire \u_ppwm/u_mem/_0062_ ;
 wire \u_ppwm/u_mem/_0063_ ;
 wire \u_ppwm/u_mem/_0064_ ;
 wire \u_ppwm/u_mem/_0065_ ;
 wire \u_ppwm/u_mem/_0066_ ;
 wire \u_ppwm/u_mem/_0067_ ;
 wire \u_ppwm/u_mem/_0068_ ;
 wire \u_ppwm/u_mem/_0069_ ;
 wire \u_ppwm/u_mem/_0070_ ;
 wire \u_ppwm/u_mem/_0071_ ;
 wire \u_ppwm/u_mem/_0072_ ;
 wire \u_ppwm/u_mem/_0073_ ;
 wire \u_ppwm/u_mem/_0074_ ;
 wire \u_ppwm/u_mem/_0075_ ;
 wire \u_ppwm/u_mem/_0076_ ;
 wire \u_ppwm/u_mem/_0077_ ;
 wire \u_ppwm/u_mem/_0078_ ;
 wire \u_ppwm/u_mem/_0079_ ;
 wire \u_ppwm/u_mem/_0080_ ;
 wire \u_ppwm/u_mem/_0081_ ;
 wire \u_ppwm/u_mem/_0082_ ;
 wire \u_ppwm/u_mem/_0083_ ;
 wire \u_ppwm/u_mem/_0084_ ;
 wire \u_ppwm/u_mem/_0085_ ;
 wire \u_ppwm/u_mem/_0086_ ;
 wire \u_ppwm/u_mem/_0087_ ;
 wire \u_ppwm/u_mem/_0088_ ;
 wire \u_ppwm/u_mem/_0089_ ;
 wire \u_ppwm/u_mem/_0090_ ;
 wire \u_ppwm/u_mem/_0091_ ;
 wire \u_ppwm/u_mem/_0092_ ;
 wire \u_ppwm/u_mem/_0093_ ;
 wire \u_ppwm/u_mem/_0094_ ;
 wire \u_ppwm/u_mem/_0095_ ;
 wire \u_ppwm/u_mem/_0096_ ;
 wire \u_ppwm/u_mem/_0097_ ;
 wire \u_ppwm/u_mem/_0098_ ;
 wire \u_ppwm/u_mem/_0099_ ;
 wire \u_ppwm/u_mem/_0100_ ;
 wire \u_ppwm/u_mem/_0101_ ;
 wire \u_ppwm/u_mem/_0102_ ;
 wire \u_ppwm/u_mem/_0103_ ;
 wire \u_ppwm/u_mem/_0104_ ;
 wire \u_ppwm/u_mem/_0105_ ;
 wire \u_ppwm/u_mem/_0106_ ;
 wire \u_ppwm/u_mem/_0107_ ;
 wire \u_ppwm/u_mem/_0108_ ;
 wire \u_ppwm/u_mem/_0109_ ;
 wire \u_ppwm/u_mem/_0110_ ;
 wire \u_ppwm/u_mem/_0111_ ;
 wire \u_ppwm/u_mem/_0112_ ;
 wire \u_ppwm/u_mem/_0113_ ;
 wire \u_ppwm/u_mem/_0114_ ;
 wire \u_ppwm/u_mem/_0115_ ;
 wire \u_ppwm/u_mem/_0116_ ;
 wire \u_ppwm/u_mem/_0117_ ;
 wire \u_ppwm/u_mem/_0118_ ;
 wire \u_ppwm/u_mem/_0119_ ;
 wire \u_ppwm/u_mem/_0120_ ;
 wire \u_ppwm/u_mem/_0121_ ;
 wire \u_ppwm/u_mem/_0122_ ;
 wire \u_ppwm/u_mem/_0123_ ;
 wire \u_ppwm/u_mem/_0124_ ;
 wire \u_ppwm/u_mem/_0125_ ;
 wire \u_ppwm/u_mem/_0126_ ;
 wire \u_ppwm/u_mem/_0127_ ;
 wire \u_ppwm/u_mem/_0128_ ;
 wire \u_ppwm/u_mem/_0129_ ;
 wire \u_ppwm/u_mem/_0130_ ;
 wire \u_ppwm/u_mem/_0131_ ;
 wire \u_ppwm/u_mem/_0132_ ;
 wire \u_ppwm/u_mem/_0133_ ;
 wire \u_ppwm/u_mem/_0134_ ;
 wire \u_ppwm/u_mem/_0135_ ;
 wire \u_ppwm/u_mem/_0136_ ;
 wire \u_ppwm/u_mem/_0137_ ;
 wire \u_ppwm/u_mem/_0138_ ;
 wire \u_ppwm/u_mem/_0139_ ;
 wire \u_ppwm/u_mem/_0140_ ;
 wire \u_ppwm/u_mem/_0141_ ;
 wire \u_ppwm/u_mem/_0142_ ;
 wire \u_ppwm/u_mem/_0143_ ;
 wire \u_ppwm/u_mem/_0144_ ;
 wire \u_ppwm/u_mem/_0145_ ;
 wire \u_ppwm/u_mem/_0146_ ;
 wire \u_ppwm/u_mem/_0147_ ;
 wire \u_ppwm/u_mem/_0148_ ;
 wire \u_ppwm/u_mem/_0149_ ;
 wire \u_ppwm/u_mem/_0150_ ;
 wire \u_ppwm/u_mem/_0151_ ;
 wire \u_ppwm/u_mem/_0152_ ;
 wire \u_ppwm/u_mem/_0153_ ;
 wire \u_ppwm/u_mem/_0154_ ;
 wire \u_ppwm/u_mem/_0155_ ;
 wire \u_ppwm/u_mem/_0156_ ;
 wire \u_ppwm/u_mem/_0157_ ;
 wire \u_ppwm/u_mem/_0158_ ;
 wire \u_ppwm/u_mem/_0159_ ;
 wire \u_ppwm/u_mem/_0160_ ;
 wire \u_ppwm/u_mem/_0161_ ;
 wire \u_ppwm/u_mem/_0162_ ;
 wire \u_ppwm/u_mem/_0163_ ;
 wire \u_ppwm/u_mem/_0164_ ;
 wire \u_ppwm/u_mem/_0165_ ;
 wire \u_ppwm/u_mem/_0166_ ;
 wire \u_ppwm/u_mem/_0167_ ;
 wire \u_ppwm/u_mem/_0168_ ;
 wire \u_ppwm/u_mem/_0169_ ;
 wire \u_ppwm/u_mem/_0170_ ;
 wire \u_ppwm/u_mem/_0171_ ;
 wire \u_ppwm/u_mem/_0172_ ;
 wire \u_ppwm/u_mem/_0173_ ;
 wire \u_ppwm/u_mem/_0174_ ;
 wire \u_ppwm/u_mem/_0175_ ;
 wire \u_ppwm/u_mem/_0176_ ;
 wire \u_ppwm/u_mem/_0177_ ;
 wire \u_ppwm/u_mem/_0178_ ;
 wire \u_ppwm/u_mem/_0179_ ;
 wire \u_ppwm/u_mem/_0180_ ;
 wire \u_ppwm/u_mem/_0181_ ;
 wire \u_ppwm/u_mem/_0182_ ;
 wire \u_ppwm/u_mem/_0183_ ;
 wire \u_ppwm/u_mem/_0184_ ;
 wire \u_ppwm/u_mem/_0185_ ;
 wire \u_ppwm/u_mem/_0186_ ;
 wire \u_ppwm/u_mem/_0187_ ;
 wire \u_ppwm/u_mem/_0188_ ;
 wire \u_ppwm/u_mem/_0189_ ;
 wire \u_ppwm/u_mem/_0190_ ;
 wire \u_ppwm/u_mem/_0191_ ;
 wire \u_ppwm/u_mem/_0192_ ;
 wire \u_ppwm/u_mem/_0193_ ;
 wire \u_ppwm/u_mem/_0194_ ;
 wire \u_ppwm/u_mem/_0195_ ;
 wire \u_ppwm/u_mem/_0196_ ;
 wire \u_ppwm/u_mem/_0197_ ;
 wire \u_ppwm/u_mem/_0198_ ;
 wire \u_ppwm/u_mem/_0199_ ;
 wire \u_ppwm/u_mem/_0200_ ;
 wire \u_ppwm/u_mem/_0201_ ;
 wire \u_ppwm/u_mem/_0202_ ;
 wire \u_ppwm/u_mem/_0203_ ;
 wire \u_ppwm/u_mem/_0204_ ;
 wire \u_ppwm/u_mem/_0205_ ;
 wire \u_ppwm/u_mem/_0206_ ;
 wire \u_ppwm/u_mem/_0207_ ;
 wire \u_ppwm/u_mem/_0208_ ;
 wire \u_ppwm/u_mem/_0209_ ;
 wire \u_ppwm/u_mem/_0210_ ;
 wire \u_ppwm/u_mem/_0211_ ;
 wire \u_ppwm/u_mem/_0212_ ;
 wire \u_ppwm/u_mem/_0213_ ;
 wire \u_ppwm/u_mem/_0214_ ;
 wire \u_ppwm/u_mem/_0215_ ;
 wire \u_ppwm/u_mem/_0216_ ;
 wire \u_ppwm/u_mem/_0217_ ;
 wire \u_ppwm/u_mem/_0218_ ;
 wire \u_ppwm/u_mem/_0219_ ;
 wire \u_ppwm/u_mem/_0220_ ;
 wire \u_ppwm/u_mem/_0221_ ;
 wire \u_ppwm/u_mem/_0222_ ;
 wire \u_ppwm/u_mem/_0223_ ;
 wire \u_ppwm/u_mem/_0224_ ;
 wire \u_ppwm/u_mem/_0225_ ;
 wire \u_ppwm/u_mem/_0226_ ;
 wire \u_ppwm/u_mem/_0227_ ;
 wire \u_ppwm/u_mem/_0228_ ;
 wire \u_ppwm/u_mem/_0229_ ;
 wire \u_ppwm/u_mem/_0230_ ;
 wire \u_ppwm/u_mem/_0231_ ;
 wire \u_ppwm/u_mem/_0232_ ;
 wire \u_ppwm/u_mem/_0233_ ;
 wire \u_ppwm/u_mem/_0234_ ;
 wire \u_ppwm/u_mem/_0235_ ;
 wire \u_ppwm/u_mem/_0236_ ;
 wire \u_ppwm/u_mem/_0237_ ;
 wire \u_ppwm/u_mem/_0238_ ;
 wire \u_ppwm/u_mem/_0239_ ;
 wire \u_ppwm/u_mem/_0240_ ;
 wire \u_ppwm/u_mem/_0241_ ;
 wire \u_ppwm/u_mem/_0242_ ;
 wire \u_ppwm/u_mem/_0243_ ;
 wire \u_ppwm/u_mem/_0244_ ;
 wire \u_ppwm/u_mem/_0245_ ;
 wire \u_ppwm/u_mem/_0246_ ;
 wire \u_ppwm/u_mem/_0247_ ;
 wire \u_ppwm/u_mem/_0248_ ;
 wire \u_ppwm/u_mem/_0249_ ;
 wire \u_ppwm/u_mem/_0250_ ;
 wire \u_ppwm/u_mem/_0251_ ;
 wire \u_ppwm/u_mem/_0252_ ;
 wire \u_ppwm/u_mem/_0253_ ;
 wire \u_ppwm/u_mem/_0254_ ;
 wire \u_ppwm/u_mem/_0255_ ;
 wire \u_ppwm/u_mem/_0256_ ;
 wire \u_ppwm/u_mem/_0257_ ;
 wire \u_ppwm/u_mem/_0258_ ;
 wire \u_ppwm/u_mem/_0259_ ;
 wire \u_ppwm/u_mem/_0260_ ;
 wire \u_ppwm/u_mem/_0261_ ;
 wire \u_ppwm/u_mem/_0262_ ;
 wire \u_ppwm/u_mem/_0263_ ;
 wire \u_ppwm/u_mem/_0264_ ;
 wire \u_ppwm/u_mem/_0265_ ;
 wire \u_ppwm/u_mem/_0266_ ;
 wire \u_ppwm/u_mem/_0267_ ;
 wire \u_ppwm/u_mem/_0268_ ;
 wire \u_ppwm/u_mem/_0269_ ;
 wire \u_ppwm/u_mem/_0270_ ;
 wire \u_ppwm/u_mem/_0271_ ;
 wire \u_ppwm/u_mem/_0272_ ;
 wire \u_ppwm/u_mem/_0273_ ;
 wire \u_ppwm/u_mem/_0274_ ;
 wire \u_ppwm/u_mem/_0275_ ;
 wire \u_ppwm/u_mem/_0276_ ;
 wire \u_ppwm/u_mem/_0277_ ;
 wire \u_ppwm/u_mem/_0278_ ;
 wire \u_ppwm/u_mem/_0279_ ;
 wire \u_ppwm/u_mem/_0280_ ;
 wire \u_ppwm/u_mem/_0281_ ;
 wire \u_ppwm/u_mem/_0282_ ;
 wire \u_ppwm/u_mem/_0283_ ;
 wire \u_ppwm/u_mem/_0284_ ;
 wire \u_ppwm/u_mem/_0285_ ;
 wire \u_ppwm/u_mem/_0286_ ;
 wire \u_ppwm/u_mem/_0287_ ;
 wire \u_ppwm/u_mem/_0288_ ;
 wire \u_ppwm/u_mem/_0289_ ;
 wire \u_ppwm/u_mem/_0290_ ;
 wire \u_ppwm/u_mem/_0291_ ;
 wire \u_ppwm/u_mem/_0292_ ;
 wire \u_ppwm/u_mem/_0293_ ;
 wire \u_ppwm/u_mem/_0294_ ;
 wire \u_ppwm/u_mem/_0295_ ;
 wire \u_ppwm/u_mem/_0296_ ;
 wire \u_ppwm/u_mem/_0297_ ;
 wire \u_ppwm/u_mem/_0298_ ;
 wire \u_ppwm/u_mem/_0299_ ;
 wire \u_ppwm/u_mem/_0300_ ;
 wire \u_ppwm/u_mem/_0301_ ;
 wire \u_ppwm/u_mem/_0302_ ;
 wire \u_ppwm/u_mem/_0303_ ;
 wire \u_ppwm/u_mem/_0304_ ;
 wire \u_ppwm/u_mem/_0305_ ;
 wire \u_ppwm/u_mem/_0306_ ;
 wire \u_ppwm/u_mem/_0307_ ;
 wire \u_ppwm/u_mem/_0308_ ;
 wire \u_ppwm/u_mem/_0309_ ;
 wire \u_ppwm/u_mem/_0310_ ;
 wire \u_ppwm/u_mem/_0311_ ;
 wire \u_ppwm/u_mem/_0312_ ;
 wire \u_ppwm/u_mem/_0313_ ;
 wire \u_ppwm/u_mem/_0314_ ;
 wire \u_ppwm/u_mem/_0315_ ;
 wire \u_ppwm/u_mem/_0316_ ;
 wire \u_ppwm/u_mem/_0317_ ;
 wire \u_ppwm/u_mem/_0318_ ;
 wire \u_ppwm/u_mem/_0319_ ;
 wire \u_ppwm/u_mem/_0320_ ;
 wire \u_ppwm/u_mem/_0321_ ;
 wire \u_ppwm/u_mem/_0322_ ;
 wire \u_ppwm/u_mem/_0323_ ;
 wire \u_ppwm/u_mem/_0324_ ;
 wire \u_ppwm/u_mem/_0325_ ;
 wire \u_ppwm/u_mem/_0326_ ;
 wire \u_ppwm/u_mem/_0327_ ;
 wire \u_ppwm/u_mem/_0328_ ;
 wire \u_ppwm/u_mem/_0329_ ;
 wire \u_ppwm/u_mem/_0330_ ;
 wire \u_ppwm/u_mem/_0331_ ;
 wire \u_ppwm/u_mem/_0332_ ;
 wire \u_ppwm/u_mem/_0333_ ;
 wire \u_ppwm/u_mem/_0334_ ;
 wire \u_ppwm/u_mem/_0335_ ;
 wire \u_ppwm/u_mem/_0336_ ;
 wire \u_ppwm/u_mem/_0337_ ;
 wire \u_ppwm/u_mem/_0338_ ;
 wire \u_ppwm/u_mem/_0339_ ;
 wire \u_ppwm/u_mem/_0340_ ;
 wire \u_ppwm/u_mem/_0341_ ;
 wire \u_ppwm/u_mem/_0342_ ;
 wire \u_ppwm/u_mem/_0343_ ;
 wire \u_ppwm/u_mem/_0344_ ;
 wire \u_ppwm/u_mem/_0345_ ;
 wire \u_ppwm/u_mem/_0346_ ;
 wire \u_ppwm/u_mem/_0347_ ;
 wire \u_ppwm/u_mem/_0348_ ;
 wire \u_ppwm/u_mem/_0349_ ;
 wire \u_ppwm/u_mem/_0350_ ;
 wire \u_ppwm/u_mem/_0351_ ;
 wire \u_ppwm/u_mem/_0352_ ;
 wire \u_ppwm/u_mem/_0353_ ;
 wire \u_ppwm/u_mem/_0354_ ;
 wire \u_ppwm/u_mem/_0355_ ;
 wire \u_ppwm/u_mem/_0356_ ;
 wire \u_ppwm/u_mem/_0357_ ;
 wire \u_ppwm/u_mem/_0358_ ;
 wire \u_ppwm/u_mem/_0359_ ;
 wire \u_ppwm/u_mem/_0360_ ;
 wire \u_ppwm/u_mem/_0361_ ;
 wire \u_ppwm/u_mem/_0362_ ;
 wire \u_ppwm/u_mem/_0363_ ;
 wire \u_ppwm/u_mem/_0364_ ;
 wire \u_ppwm/u_mem/_0365_ ;
 wire \u_ppwm/u_mem/_0366_ ;
 wire \u_ppwm/u_mem/_0367_ ;
 wire \u_ppwm/u_mem/_0368_ ;
 wire \u_ppwm/u_mem/_0369_ ;
 wire \u_ppwm/u_mem/_0370_ ;
 wire \u_ppwm/u_mem/_0371_ ;
 wire \u_ppwm/u_mem/_0372_ ;
 wire \u_ppwm/u_mem/_0373_ ;
 wire \u_ppwm/u_mem/_0374_ ;
 wire \u_ppwm/u_mem/_0375_ ;
 wire \u_ppwm/u_mem/_0376_ ;
 wire \u_ppwm/u_mem/_0377_ ;
 wire \u_ppwm/u_mem/_0378_ ;
 wire \u_ppwm/u_mem/_0379_ ;
 wire \u_ppwm/u_mem/_0380_ ;
 wire \u_ppwm/u_mem/_0381_ ;
 wire \u_ppwm/u_mem/_0382_ ;
 wire \u_ppwm/u_mem/_0383_ ;
 wire \u_ppwm/u_mem/_0384_ ;
 wire \u_ppwm/u_mem/_0385_ ;
 wire \u_ppwm/u_mem/_0386_ ;
 wire \u_ppwm/u_mem/_0387_ ;
 wire \u_ppwm/u_mem/_0388_ ;
 wire \u_ppwm/u_mem/_0389_ ;
 wire \u_ppwm/u_mem/_0390_ ;
 wire \u_ppwm/u_mem/_0391_ ;
 wire \u_ppwm/u_mem/_0392_ ;
 wire \u_ppwm/u_mem/_0393_ ;
 wire \u_ppwm/u_mem/_0394_ ;
 wire \u_ppwm/u_mem/_0395_ ;
 wire \u_ppwm/u_mem/_0396_ ;
 wire \u_ppwm/u_mem/_0397_ ;
 wire \u_ppwm/u_mem/_0398_ ;
 wire \u_ppwm/u_mem/_0399_ ;
 wire \u_ppwm/u_mem/_0400_ ;
 wire \u_ppwm/u_mem/_0401_ ;
 wire \u_ppwm/u_mem/_0402_ ;
 wire \u_ppwm/u_mem/_0403_ ;
 wire \u_ppwm/u_mem/_0404_ ;
 wire \u_ppwm/u_mem/_0405_ ;
 wire \u_ppwm/u_mem/_0406_ ;
 wire \u_ppwm/u_mem/_0407_ ;
 wire \u_ppwm/u_mem/_0408_ ;
 wire \u_ppwm/u_mem/_0409_ ;
 wire \u_ppwm/u_mem/_0410_ ;
 wire \u_ppwm/u_mem/_0411_ ;
 wire \u_ppwm/u_mem/_0412_ ;
 wire \u_ppwm/u_mem/_0413_ ;
 wire \u_ppwm/u_mem/_0414_ ;
 wire \u_ppwm/u_mem/_0415_ ;
 wire \u_ppwm/u_mem/_0416_ ;
 wire \u_ppwm/u_mem/_0417_ ;
 wire \u_ppwm/u_mem/_0418_ ;
 wire \u_ppwm/u_mem/_0419_ ;
 wire \u_ppwm/u_mem/_0420_ ;
 wire \u_ppwm/u_mem/_0421_ ;
 wire \u_ppwm/u_mem/_0422_ ;
 wire \u_ppwm/u_mem/_0423_ ;
 wire \u_ppwm/u_mem/_0424_ ;
 wire \u_ppwm/u_mem/_0425_ ;
 wire \u_ppwm/u_mem/_0426_ ;
 wire \u_ppwm/u_mem/_0427_ ;
 wire \u_ppwm/u_mem/_0428_ ;
 wire \u_ppwm/u_mem/_0429_ ;
 wire \u_ppwm/u_mem/_0430_ ;
 wire \u_ppwm/u_mem/_0431_ ;
 wire \u_ppwm/u_mem/_0432_ ;
 wire \u_ppwm/u_mem/_0433_ ;
 wire \u_ppwm/u_mem/_0434_ ;
 wire \u_ppwm/u_mem/_0435_ ;
 wire \u_ppwm/u_mem/_0436_ ;
 wire \u_ppwm/u_mem/_0437_ ;
 wire \u_ppwm/u_mem/_0438_ ;
 wire \u_ppwm/u_mem/_0439_ ;
 wire \u_ppwm/u_mem/_0440_ ;
 wire \u_ppwm/u_mem/_0441_ ;
 wire \u_ppwm/u_mem/_0442_ ;
 wire \u_ppwm/u_mem/_0443_ ;
 wire \u_ppwm/u_mem/_0444_ ;
 wire \u_ppwm/u_mem/_0445_ ;
 wire \u_ppwm/u_mem/_0446_ ;
 wire \u_ppwm/u_mem/_0447_ ;
 wire \u_ppwm/u_mem/_0448_ ;
 wire \u_ppwm/u_mem/_0449_ ;
 wire \u_ppwm/u_mem/_0450_ ;
 wire \u_ppwm/u_mem/_0451_ ;
 wire \u_ppwm/u_mem/_0452_ ;
 wire \u_ppwm/u_mem/_0453_ ;
 wire \u_ppwm/u_mem/_0454_ ;
 wire \u_ppwm/u_mem/_0455_ ;
 wire \u_ppwm/u_mem/_0456_ ;
 wire \u_ppwm/u_mem/_0457_ ;
 wire \u_ppwm/u_mem/_0458_ ;
 wire \u_ppwm/u_mem/_0459_ ;
 wire \u_ppwm/u_mem/_0460_ ;
 wire \u_ppwm/u_mem/_0461_ ;
 wire \u_ppwm/u_mem/_0462_ ;
 wire \u_ppwm/u_mem/_0463_ ;
 wire \u_ppwm/u_mem/_0464_ ;
 wire \u_ppwm/u_mem/_0465_ ;
 wire \u_ppwm/u_mem/_0466_ ;
 wire \u_ppwm/u_mem/_0467_ ;
 wire \u_ppwm/u_mem/_0468_ ;
 wire \u_ppwm/u_mem/_0469_ ;
 wire \u_ppwm/u_mem/_0470_ ;
 wire \u_ppwm/u_mem/_0471_ ;
 wire \u_ppwm/u_mem/_0472_ ;
 wire \u_ppwm/u_mem/_0473_ ;
 wire \u_ppwm/u_mem/_0474_ ;
 wire \u_ppwm/u_mem/_0475_ ;
 wire \u_ppwm/u_mem/_0476_ ;
 wire \u_ppwm/u_mem/_0477_ ;
 wire \u_ppwm/u_mem/_0478_ ;
 wire \u_ppwm/u_mem/_0479_ ;
 wire \u_ppwm/u_mem/_0480_ ;
 wire \u_ppwm/u_mem/_0481_ ;
 wire \u_ppwm/u_mem/_0482_ ;
 wire \u_ppwm/u_mem/_0483_ ;
 wire \u_ppwm/u_mem/_0484_ ;
 wire \u_ppwm/u_mem/_0485_ ;
 wire \u_ppwm/u_mem/_0486_ ;
 wire \u_ppwm/u_mem/_0487_ ;
 wire \u_ppwm/u_mem/_0488_ ;
 wire \u_ppwm/u_mem/_0489_ ;
 wire \u_ppwm/u_mem/_0490_ ;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire \u_ppwm/u_mem/bit_count[0] ;
 wire \u_ppwm/u_mem/bit_count[1] ;
 wire \u_ppwm/u_mem/bit_count[2] ;
 wire \u_ppwm/u_mem/bit_count[3] ;
 wire \u_ppwm/u_mem/bit_count[4] ;
 wire \u_ppwm/u_mem/bit_count[5] ;
 wire \u_ppwm/u_mem/bit_count[6] ;
 wire \u_ppwm/u_mem/memory[0] ;
 wire \u_ppwm/u_mem/memory[100] ;
 wire \u_ppwm/u_mem/memory[101] ;
 wire \u_ppwm/u_mem/memory[102] ;
 wire \u_ppwm/u_mem/memory[103] ;
 wire \u_ppwm/u_mem/memory[104] ;
 wire \u_ppwm/u_mem/memory[105] ;
 wire \u_ppwm/u_mem/memory[106] ;
 wire \u_ppwm/u_mem/memory[107] ;
 wire \u_ppwm/u_mem/memory[10] ;
 wire \u_ppwm/u_mem/memory[11] ;
 wire \u_ppwm/u_mem/memory[12] ;
 wire \u_ppwm/u_mem/memory[13] ;
 wire \u_ppwm/u_mem/memory[14] ;
 wire \u_ppwm/u_mem/memory[15] ;
 wire \u_ppwm/u_mem/memory[16] ;
 wire \u_ppwm/u_mem/memory[17] ;
 wire \u_ppwm/u_mem/memory[18] ;
 wire \u_ppwm/u_mem/memory[19] ;
 wire \u_ppwm/u_mem/memory[1] ;
 wire \u_ppwm/u_mem/memory[20] ;
 wire \u_ppwm/u_mem/memory[21] ;
 wire \u_ppwm/u_mem/memory[22] ;
 wire \u_ppwm/u_mem/memory[23] ;
 wire \u_ppwm/u_mem/memory[24] ;
 wire \u_ppwm/u_mem/memory[25] ;
 wire \u_ppwm/u_mem/memory[26] ;
 wire \u_ppwm/u_mem/memory[27] ;
 wire \u_ppwm/u_mem/memory[28] ;
 wire \u_ppwm/u_mem/memory[29] ;
 wire \u_ppwm/u_mem/memory[2] ;
 wire \u_ppwm/u_mem/memory[30] ;
 wire \u_ppwm/u_mem/memory[31] ;
 wire \u_ppwm/u_mem/memory[32] ;
 wire \u_ppwm/u_mem/memory[33] ;
 wire \u_ppwm/u_mem/memory[34] ;
 wire \u_ppwm/u_mem/memory[35] ;
 wire \u_ppwm/u_mem/memory[36] ;
 wire \u_ppwm/u_mem/memory[37] ;
 wire \u_ppwm/u_mem/memory[38] ;
 wire \u_ppwm/u_mem/memory[39] ;
 wire \u_ppwm/u_mem/memory[3] ;
 wire \u_ppwm/u_mem/memory[40] ;
 wire \u_ppwm/u_mem/memory[41] ;
 wire \u_ppwm/u_mem/memory[42] ;
 wire \u_ppwm/u_mem/memory[43] ;
 wire \u_ppwm/u_mem/memory[44] ;
 wire \u_ppwm/u_mem/memory[45] ;
 wire \u_ppwm/u_mem/memory[46] ;
 wire \u_ppwm/u_mem/memory[47] ;
 wire \u_ppwm/u_mem/memory[48] ;
 wire \u_ppwm/u_mem/memory[49] ;
 wire \u_ppwm/u_mem/memory[4] ;
 wire \u_ppwm/u_mem/memory[50] ;
 wire \u_ppwm/u_mem/memory[51] ;
 wire \u_ppwm/u_mem/memory[52] ;
 wire \u_ppwm/u_mem/memory[53] ;
 wire \u_ppwm/u_mem/memory[54] ;
 wire \u_ppwm/u_mem/memory[55] ;
 wire \u_ppwm/u_mem/memory[56] ;
 wire \u_ppwm/u_mem/memory[57] ;
 wire \u_ppwm/u_mem/memory[58] ;
 wire \u_ppwm/u_mem/memory[59] ;
 wire \u_ppwm/u_mem/memory[5] ;
 wire \u_ppwm/u_mem/memory[60] ;
 wire \u_ppwm/u_mem/memory[61] ;
 wire \u_ppwm/u_mem/memory[62] ;
 wire \u_ppwm/u_mem/memory[63] ;
 wire \u_ppwm/u_mem/memory[64] ;
 wire \u_ppwm/u_mem/memory[65] ;
 wire \u_ppwm/u_mem/memory[66] ;
 wire \u_ppwm/u_mem/memory[67] ;
 wire \u_ppwm/u_mem/memory[68] ;
 wire \u_ppwm/u_mem/memory[69] ;
 wire \u_ppwm/u_mem/memory[6] ;
 wire \u_ppwm/u_mem/memory[70] ;
 wire \u_ppwm/u_mem/memory[71] ;
 wire \u_ppwm/u_mem/memory[72] ;
 wire \u_ppwm/u_mem/memory[73] ;
 wire \u_ppwm/u_mem/memory[74] ;
 wire \u_ppwm/u_mem/memory[75] ;
 wire \u_ppwm/u_mem/memory[76] ;
 wire \u_ppwm/u_mem/memory[77] ;
 wire \u_ppwm/u_mem/memory[78] ;
 wire \u_ppwm/u_mem/memory[79] ;
 wire \u_ppwm/u_mem/memory[7] ;
 wire \u_ppwm/u_mem/memory[80] ;
 wire \u_ppwm/u_mem/memory[81] ;
 wire \u_ppwm/u_mem/memory[82] ;
 wire \u_ppwm/u_mem/memory[83] ;
 wire \u_ppwm/u_mem/memory[84] ;
 wire \u_ppwm/u_mem/memory[85] ;
 wire \u_ppwm/u_mem/memory[86] ;
 wire \u_ppwm/u_mem/memory[87] ;
 wire \u_ppwm/u_mem/memory[88] ;
 wire \u_ppwm/u_mem/memory[89] ;
 wire \u_ppwm/u_mem/memory[8] ;
 wire \u_ppwm/u_mem/memory[90] ;
 wire \u_ppwm/u_mem/memory[91] ;
 wire \u_ppwm/u_mem/memory[92] ;
 wire \u_ppwm/u_mem/memory[93] ;
 wire \u_ppwm/u_mem/memory[94] ;
 wire \u_ppwm/u_mem/memory[95] ;
 wire \u_ppwm/u_mem/memory[96] ;
 wire \u_ppwm/u_mem/memory[97] ;
 wire \u_ppwm/u_mem/memory[98] ;
 wire \u_ppwm/u_mem/memory[99] ;
 wire \u_ppwm/u_mem/memory[9] ;
 wire \u_ppwm/u_mem/state_q[0] ;
 wire \u_ppwm/u_mem/state_q[2] ;
 wire \u_ppwm/u_pwm/_000_ ;
 wire \u_ppwm/u_pwm/_001_ ;
 wire \u_ppwm/u_pwm/_002_ ;
 wire \u_ppwm/u_pwm/_003_ ;
 wire \u_ppwm/u_pwm/_004_ ;
 wire \u_ppwm/u_pwm/_005_ ;
 wire \u_ppwm/u_pwm/_006_ ;
 wire \u_ppwm/u_pwm/_007_ ;
 wire \u_ppwm/u_pwm/_008_ ;
 wire \u_ppwm/u_pwm/_009_ ;
 wire \u_ppwm/u_pwm/_010_ ;
 wire \u_ppwm/u_pwm/_011_ ;
 wire \u_ppwm/u_pwm/_012_ ;
 wire \u_ppwm/u_pwm/_013_ ;
 wire \u_ppwm/u_pwm/_014_ ;
 wire \u_ppwm/u_pwm/_015_ ;
 wire \u_ppwm/u_pwm/_016_ ;
 wire \u_ppwm/u_pwm/_017_ ;
 wire \u_ppwm/u_pwm/_018_ ;
 wire \u_ppwm/u_pwm/_019_ ;
 wire \u_ppwm/u_pwm/_020_ ;
 wire \u_ppwm/u_pwm/_021_ ;
 wire \u_ppwm/u_pwm/_022_ ;
 wire \u_ppwm/u_pwm/_023_ ;
 wire \u_ppwm/u_pwm/_024_ ;
 wire \u_ppwm/u_pwm/_025_ ;
 wire \u_ppwm/u_pwm/_026_ ;
 wire \u_ppwm/u_pwm/_027_ ;
 wire \u_ppwm/u_pwm/_028_ ;
 wire \u_ppwm/u_pwm/_029_ ;
 wire \u_ppwm/u_pwm/_030_ ;
 wire \u_ppwm/u_pwm/_031_ ;
 wire \u_ppwm/u_pwm/_032_ ;
 wire \u_ppwm/u_pwm/_033_ ;
 wire \u_ppwm/u_pwm/_034_ ;
 wire \u_ppwm/u_pwm/_035_ ;
 wire \u_ppwm/u_pwm/_036_ ;
 wire \u_ppwm/u_pwm/_037_ ;
 wire \u_ppwm/u_pwm/_038_ ;
 wire \u_ppwm/u_pwm/_039_ ;
 wire \u_ppwm/u_pwm/_040_ ;
 wire \u_ppwm/u_pwm/_041_ ;
 wire \u_ppwm/u_pwm/_042_ ;
 wire \u_ppwm/u_pwm/_043_ ;
 wire \u_ppwm/u_pwm/_044_ ;
 wire \u_ppwm/u_pwm/_045_ ;
 wire \u_ppwm/u_pwm/_046_ ;
 wire \u_ppwm/u_pwm/_047_ ;
 wire \u_ppwm/u_pwm/_048_ ;
 wire \u_ppwm/u_pwm/_049_ ;
 wire \u_ppwm/u_pwm/_050_ ;
 wire \u_ppwm/u_pwm/_051_ ;
 wire \u_ppwm/u_pwm/_052_ ;
 wire \u_ppwm/u_pwm/_053_ ;
 wire \u_ppwm/u_pwm/_054_ ;
 wire \u_ppwm/u_pwm/_055_ ;
 wire \u_ppwm/u_pwm/_056_ ;
 wire \u_ppwm/u_pwm/_057_ ;
 wire \u_ppwm/u_pwm/_058_ ;
 wire \u_ppwm/u_pwm/_059_ ;
 wire \u_ppwm/u_pwm/_060_ ;
 wire \u_ppwm/u_pwm/_061_ ;
 wire \u_ppwm/u_pwm/_062_ ;
 wire \u_ppwm/u_pwm/_063_ ;
 wire \u_ppwm/u_pwm/_064_ ;
 wire \u_ppwm/u_pwm/_065_ ;
 wire \u_ppwm/u_pwm/_066_ ;
 wire \u_ppwm/u_pwm/_067_ ;
 wire \u_ppwm/u_pwm/_068_ ;
 wire \u_ppwm/u_pwm/_069_ ;
 wire \u_ppwm/u_pwm/_070_ ;
 wire \u_ppwm/u_pwm/_071_ ;
 wire \u_ppwm/u_pwm/_072_ ;
 wire \u_ppwm/u_pwm/_073_ ;
 wire \u_ppwm/u_pwm/_074_ ;
 wire \u_ppwm/u_pwm/_075_ ;
 wire \u_ppwm/u_pwm/_076_ ;
 wire \u_ppwm/u_pwm/_077_ ;
 wire \u_ppwm/u_pwm/_078_ ;
 wire \u_ppwm/u_pwm/_079_ ;
 wire \u_ppwm/u_pwm/_080_ ;
 wire \u_ppwm/u_pwm/_081_ ;
 wire \u_ppwm/u_pwm/_082_ ;
 wire \u_ppwm/u_pwm/_083_ ;
 wire \u_ppwm/u_pwm/_084_ ;
 wire \u_ppwm/u_pwm/_085_ ;
 wire \u_ppwm/u_pwm/_086_ ;
 wire \u_ppwm/u_pwm/_087_ ;
 wire \u_ppwm/u_pwm/_088_ ;
 wire \u_ppwm/u_pwm/_089_ ;
 wire \u_ppwm/u_pwm/_090_ ;
 wire \u_ppwm/u_pwm/_091_ ;
 wire \u_ppwm/u_pwm/_092_ ;
 wire \u_ppwm/u_pwm/_093_ ;
 wire \u_ppwm/u_pwm/_094_ ;
 wire \u_ppwm/u_pwm/_095_ ;
 wire \u_ppwm/u_pwm/_096_ ;
 wire \u_ppwm/u_pwm/_097_ ;
 wire \u_ppwm/u_pwm/_098_ ;
 wire \u_ppwm/u_pwm/_099_ ;
 wire \u_ppwm/u_pwm/_100_ ;
 wire \u_ppwm/u_pwm/_101_ ;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire clknet_0_clk;
 wire \u_ppwm/u_pwm/cmp_value[0] ;
 wire \u_ppwm/u_pwm/cmp_value[1] ;
 wire \u_ppwm/u_pwm/cmp_value[2] ;
 wire \u_ppwm/u_pwm/cmp_value[3] ;
 wire \u_ppwm/u_pwm/cmp_value[4] ;
 wire \u_ppwm/u_pwm/cmp_value[5] ;
 wire \u_ppwm/u_pwm/cmp_value[6] ;
 wire \u_ppwm/u_pwm/cmp_value[7] ;
 wire \u_ppwm/u_pwm/cmp_value[8] ;
 wire \u_ppwm/u_pwm/cmp_value[9] ;
 wire \u_ppwm/u_pwm/counter[0] ;
 wire \u_ppwm/u_pwm/counter[1] ;
 wire \u_ppwm/u_pwm/counter[2] ;
 wire \u_ppwm/u_pwm/counter[3] ;
 wire \u_ppwm/u_pwm/counter[4] ;
 wire \u_ppwm/u_pwm/counter[5] ;
 wire \u_ppwm/u_pwm/counter[6] ;
 wire \u_ppwm/u_pwm/counter[7] ;
 wire \u_ppwm/u_pwm/counter[8] ;
 wire \u_ppwm/u_pwm/counter[9] ;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net1;
 wire net3;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;

 sg13g2_tielo heichips25_ppwm_4 (.L_LO(net4));
 sg13g2_tielo heichips25_ppwm_5 (.L_LO(net5));
 sg13g2_tielo heichips25_ppwm_6 (.L_LO(net6));
 sg13g2_tielo heichips25_ppwm_7 (.L_LO(net7));
 sg13g2_tielo heichips25_ppwm_8 (.L_LO(net8));
 sg13g2_tielo heichips25_ppwm_9 (.L_LO(net9));
 sg13g2_tielo heichips25_ppwm_10 (.L_LO(net10));
 sg13g2_tielo heichips25_ppwm_11 (.L_LO(net11));
 sg13g2_tielo heichips25_ppwm_12 (.L_LO(net12));
 sg13g2_tielo heichips25_ppwm_13 (.L_LO(net13));
 sg13g2_tielo heichips25_ppwm_14 (.L_LO(net14));
 sg13g2_tielo heichips25_ppwm_15 (.L_LO(net15));
 sg13g2_tielo heichips25_ppwm_16 (.L_LO(net16));
 sg13g2_tielo heichips25_ppwm_17 (.L_LO(net17));
 sg13g2_tielo heichips25_ppwm_18 (.L_LO(net18));
 sg13g2_tielo heichips25_ppwm_19 (.L_LO(net19));
 sg13g2_tielo heichips25_ppwm_20 (.L_LO(net20));
 sg13g2_tielo heichips25_ppwm_21 (.L_LO(net21));
 sg13g2_tielo heichips25_ppwm_22 (.L_LO(net22));
 sg13g2_tielo heichips25_ppwm_23 (.L_LO(net23));
 sg13g2_tielo heichips25_ppwm_24 (.L_LO(net24));
 sg13g2_tielo heichips25_ppwm_25 (.L_LO(net25));
 sg13g2_tiehi \u_ppwm/u_ex/_812__26  (.L_HI(net26));
 sg13g2_inv_2 \u_ppwm/u_ex/_415_  (.Y(\u_ppwm/u_ex/_373_ ),
    .A(\u_ppwm/u_ex/reg_value_q[7] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_416_  (.Y(\u_ppwm/u_ex/_374_ ),
    .A(net380));
 sg13g2_inv_1 \u_ppwm/u_ex/_417_  (.Y(\u_ppwm/u_ex/_375_ ),
    .A(net381));
 sg13g2_inv_1 \u_ppwm/u_ex/_418_  (.Y(\u_ppwm/u_ex/_376_ ),
    .A(net382));
 sg13g2_inv_1 \u_ppwm/u_ex/_419_  (.Y(\u_ppwm/u_ex/_377_ ),
    .A(net383));
 sg13g2_inv_2 \u_ppwm/u_ex/_420_  (.Y(\u_ppwm/u_ex/_378_ ),
    .A(net384));
 sg13g2_inv_1 \u_ppwm/u_ex/_421_  (.Y(\u_ppwm/u_ex/_379_ ),
    .A(\u_ppwm/pwm_value[9] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_422_  (.Y(\u_ppwm/u_ex/_380_ ),
    .A(net386));
 sg13g2_inv_2 \u_ppwm/u_ex/_423_  (.Y(\u_ppwm/u_ex/_381_ ),
    .A(net391));
 sg13g2_inv_1 \u_ppwm/u_ex/_424_  (.Y(\u_ppwm/u_ex/_382_ ),
    .A(net392));
 sg13g2_inv_1 \u_ppwm/u_ex/_425_  (.Y(\u_ppwm/u_ex/_383_ ),
    .A(net396));
 sg13g2_inv_1 \u_ppwm/u_ex/_426_  (.Y(\u_ppwm/u_ex/_384_ ),
    .A(net415));
 sg13g2_inv_2 \u_ppwm/u_ex/_427_  (.Y(\u_ppwm/u_ex/_385_ ),
    .A(\u_ppwm/instr[0] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_428_  (.Y(\u_ppwm/u_ex/_386_ ),
    .A(net325));
 sg13g2_inv_1 \u_ppwm/u_ex/_429_  (.Y(\u_ppwm/u_ex/_028_ ),
    .A(net336));
 sg13g2_inv_1 \u_ppwm/u_ex/_430_  (.Y(\u_ppwm/u_ex/_029_ ),
    .A(\u_ppwm/global_counter_high[16] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_431_  (.Y(\u_ppwm/u_ex/_030_ ),
    .A(\u_ppwm/global_counter_high[14] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_432_  (.Y(\u_ppwm/u_ex/_031_ ),
    .A(\u_ppwm/global_counter_high[13] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_433_  (.Y(\u_ppwm/u_ex/_032_ ),
    .A(\u_ppwm/global_counter_high[12] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_434_  (.Y(\u_ppwm/u_ex/_033_ ),
    .A(\u_ppwm/global_counter_high[9] ));
 sg13g2_inv_2 \u_ppwm/u_ex/_435_  (.Y(\u_ppwm/u_ex/_034_ ),
    .A(\u_ppwm/global_counter_high[8] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_436_  (.Y(\u_ppwm/u_ex/_035_ ),
    .A(\u_ppwm/global_counter_high[7] ));
 sg13g2_inv_2 \u_ppwm/u_ex/_437_  (.Y(\u_ppwm/u_ex/_036_ ),
    .A(\u_ppwm/global_counter_high[6] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_438_  (.Y(\u_ppwm/u_ex/_037_ ),
    .A(\u_ppwm/global_counter_high[4] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_439_  (.Y(\u_ppwm/u_ex/_038_ ),
    .A(\u_ppwm/global_counter_high[3] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_440_  (.Y(\u_ppwm/u_ex/_039_ ),
    .A(\u_ppwm/global_counter_high[2] ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_441_  (.Y(\u_ppwm/u_ex/_040_ ),
    .A(net407),
    .B(net413));
 sg13g2_nand3_1 \u_ppwm/u_ex/_442_  (.B(net406),
    .C(net412),
    .A(net402),
    .Y(\u_ppwm/u_ex/_041_ ));
 sg13g2_nand4_1 \u_ppwm/u_ex/_443_  (.B(net402),
    .C(net406),
    .A(net400),
    .Y(\u_ppwm/u_ex/_042_ ),
    .D(net413));
 sg13g2_inv_1 \u_ppwm/u_ex/_444_  (.Y(\u_ppwm/u_ex/_043_ ),
    .A(\u_ppwm/u_ex/_042_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_445_  (.A(net325),
    .B_N(net327),
    .Y(\u_ppwm/u_ex/_044_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_446_  (.Y(\u_ppwm/u_ex/_045_ ),
    .B(\u_ppwm/u_ex/_044_ ),
    .A_N(net324));
 sg13g2_or2_1 \u_ppwm/u_ex/_447_  (.X(\u_ppwm/u_ex/_046_ ),
    .B(\u_ppwm/instr[1] ),
    .A(\u_ppwm/instr[0] ));
 sg13g2_nor4_1 \u_ppwm/u_ex/_448_  (.A(\u_ppwm/instr[2] ),
    .B(net320),
    .C(\u_ppwm/u_ex/_045_ ),
    .D(\u_ppwm/u_ex/_046_ ),
    .Y(\u_ppwm/u_ex/_047_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_449_  (.Y(\u_ppwm/u_ex/_048_ ),
    .B(net377),
    .A_N(\u_ppwm/u_ex/_047_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_450_  (.B1(net427),
    .Y(\u_ppwm/u_ex/_049_ ),
    .A1(\u_ppwm/u_ex/_042_ ),
    .A2(\u_ppwm/u_ex/_048_ ));
 sg13g2_a21o_1 \u_ppwm/u_ex/_451_  (.A2(net572),
    .A1(\u_ppwm/u_ex/_028_ ),
    .B1(\u_ppwm/u_ex/_049_ ),
    .X(\u_ppwm/u_ex/_000_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_452_  (.B1(net336),
    .Y(\u_ppwm/u_ex/_050_ ),
    .A1(net572),
    .A2(net607));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_453_  (.B1(\u_ppwm/u_ex/_050_ ),
    .Y(\u_ppwm/u_ex/_051_ ),
    .A1(\u_ppwm/u_ex/_043_ ),
    .A2(\u_ppwm/u_ex/_048_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_454_  (.A(net427),
    .B(\u_ppwm/u_ex/_051_ ),
    .X(\u_ppwm/u_ex/_002_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_455_  (.Y(\u_ppwm/u_ex/_052_ ),
    .B1(\u_ppwm/u_ex/_047_ ),
    .B2(net377),
    .A2(net607),
    .A1(\u_ppwm/u_ex/_028_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_456_  (.A(net608),
    .B_N(net426),
    .Y(\u_ppwm/u_ex/_001_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_457_  (.Y(\u_ppwm/u_ex/_053_ ),
    .B(\u_ppwm/instr[1] ),
    .A_N(\u_ppwm/u_ex/cmp_flag_q ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_458_  (.B(\u_ppwm/instr[0] ),
    .C(\u_ppwm/u_ex/_053_ ),
    .A(\u_ppwm/instr[2] ),
    .Y(\u_ppwm/u_ex/_054_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_459_  (.B1(net377),
    .Y(\u_ppwm/u_ex/_055_ ),
    .A1(net327),
    .A2(\u_ppwm/u_ex/_054_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_460_  (.B1(net443),
    .Y(\u_ppwm/u_ex/_056_ ),
    .A1(\u_ppwm/u_ex/_384_ ),
    .A2(\u_ppwm/u_ex/_055_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_461_  (.A1(\u_ppwm/u_ex/_384_ ),
    .A2(\u_ppwm/u_ex/_055_ ),
    .Y(\u_ppwm/u_ex/_003_ ),
    .B1(\u_ppwm/u_ex/_056_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_462_  (.Y(\u_ppwm/u_ex/_057_ ),
    .A(\u_ppwm/u_ex/_040_ ),
    .B(\u_ppwm/u_ex/_054_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_463_  (.Y(\u_ppwm/u_ex/_058_ ),
    .A(net377),
    .B(\u_ppwm/u_ex/_057_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_464_  (.B1(\u_ppwm/u_ex/_058_ ),
    .Y(\u_ppwm/u_ex/_059_ ),
    .A1(net407),
    .A2(net415));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_465_  (.Y(\u_ppwm/u_ex/_060_ ),
    .A(net407),
    .B(net326));
 sg13g2_nand2_1 \u_ppwm/u_ex/_466_  (.Y(\u_ppwm/u_ex/_061_ ),
    .A(net415),
    .B(\u_ppwm/instr[3] ));
 sg13g2_and2_1 \u_ppwm/u_ex/_467_  (.A(\u_ppwm/u_ex/_060_ ),
    .B(\u_ppwm/u_ex/_061_ ),
    .X(\u_ppwm/u_ex/_062_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_468_  (.A(\u_ppwm/u_ex/_060_ ),
    .B(\u_ppwm/u_ex/_061_ ),
    .Y(\u_ppwm/u_ex/_063_ ));
 sg13g2_or3_1 \u_ppwm/u_ex/_469_  (.A(\u_ppwm/u_ex/_054_ ),
    .B(\u_ppwm/u_ex/_062_ ),
    .C(\u_ppwm/u_ex/_063_ ),
    .X(\u_ppwm/u_ex/_064_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_470_  (.B1(net443),
    .Y(\u_ppwm/u_ex/_065_ ),
    .A1(net377),
    .A2(net407));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_471_  (.A1(\u_ppwm/u_ex/_059_ ),
    .A2(\u_ppwm/u_ex/_064_ ),
    .Y(\u_ppwm/u_ex/_004_ ),
    .B1(\u_ppwm/u_ex/_065_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_472_  (.Y(\u_ppwm/u_ex/_066_ ),
    .B(\u_ppwm/u_ex/_040_ ),
    .A_N(net402));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_473_  (.Y(\u_ppwm/u_ex/_067_ ),
    .B(\u_ppwm/u_ex/_054_ ),
    .A_N(net402));
 sg13g2_nand3_1 \u_ppwm/u_ex/_474_  (.B(\u_ppwm/u_ex/_057_ ),
    .C(\u_ppwm/u_ex/_067_ ),
    .A(net377),
    .Y(\u_ppwm/u_ex/_068_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_475_  (.A1(net407),
    .A2(net326),
    .Y(\u_ppwm/u_ex/_069_ ),
    .B1(\u_ppwm/u_ex/_063_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_476_  (.Y(\u_ppwm/u_ex/_070_ ),
    .A(net402),
    .B(net323));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_477_  (.Y(\u_ppwm/u_ex/_071_ ),
    .A(net402),
    .B(net323));
 sg13g2_or2_1 \u_ppwm/u_ex/_478_  (.X(\u_ppwm/u_ex/_072_ ),
    .B(\u_ppwm/u_ex/_071_ ),
    .A(\u_ppwm/u_ex/_069_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_479_  (.A1(\u_ppwm/u_ex/_069_ ),
    .A2(\u_ppwm/u_ex/_071_ ),
    .Y(\u_ppwm/u_ex/_073_ ),
    .B1(\u_ppwm/u_ex/_054_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_480_  (.Y(\u_ppwm/u_ex/_074_ ),
    .B1(\u_ppwm/u_ex/_072_ ),
    .B2(\u_ppwm/u_ex/_073_ ),
    .A2(\u_ppwm/u_ex/_068_ ),
    .A1(\u_ppwm/u_ex/_066_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_481_  (.B1(net443),
    .Y(\u_ppwm/u_ex/_075_ ),
    .A1(net631),
    .A2(net402));
 sg13g2_nor2_1 \u_ppwm/u_ex/_482_  (.A(\u_ppwm/u_ex/_074_ ),
    .B(\u_ppwm/u_ex/_075_ ),
    .Y(\u_ppwm/u_ex/_005_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_483_  (.Y(\u_ppwm/u_ex/_076_ ),
    .A(net400),
    .B(net320));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_484_  (.A1(\u_ppwm/u_ex/_070_ ),
    .A2(\u_ppwm/u_ex/_072_ ),
    .Y(\u_ppwm/u_ex/_077_ ),
    .B1(\u_ppwm/u_ex/_076_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_485_  (.B(\u_ppwm/u_ex/_072_ ),
    .C(\u_ppwm/u_ex/_076_ ),
    .A(\u_ppwm/u_ex/_070_ ),
    .Y(\u_ppwm/u_ex/_078_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_486_  (.A(\u_ppwm/u_ex/_054_ ),
    .B(\u_ppwm/u_ex/_077_ ),
    .Y(\u_ppwm/u_ex/_079_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_487_  (.A(net400),
    .B_N(\u_ppwm/u_ex/_041_ ),
    .Y(\u_ppwm/u_ex/_080_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_488_  (.Y(\u_ppwm/u_ex/_081_ ),
    .A(\u_ppwm/u_ex/_042_ ),
    .B(\u_ppwm/u_ex/_054_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_489_  (.B1(net631),
    .Y(\u_ppwm/u_ex/_082_ ),
    .A1(\u_ppwm/u_ex/_080_ ),
    .A2(\u_ppwm/u_ex/_081_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_490_  (.A1(\u_ppwm/u_ex/_078_ ),
    .A2(\u_ppwm/u_ex/_079_ ),
    .Y(\u_ppwm/u_ex/_083_ ),
    .B1(\u_ppwm/u_ex/_082_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_491_  (.B1(net443),
    .Y(\u_ppwm/u_ex/_084_ ),
    .A1(net401),
    .A2(net631));
 sg13g2_nor2_1 \u_ppwm/u_ex/_492_  (.A(\u_ppwm/u_ex/_083_ ),
    .B(net632),
    .Y(\u_ppwm/u_ex/_006_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_493_  (.Y(\u_ppwm/u_ex/_085_ ),
    .B1(net198),
    .B2(\u_ppwm/u_ex/_374_ ),
    .A2(net614),
    .A1(\u_ppwm/u_ex/_373_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_494_  (.Y(\u_ppwm/u_ex/_086_ ),
    .A(net382),
    .B(\u_ppwm/u_ex/_030_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_495_  (.A(net385),
    .B_N(\u_ppwm/global_counter_high[11] ),
    .Y(\u_ppwm/u_ex/_087_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_496_  (.Y(\u_ppwm/u_ex/_088_ ),
    .B(\u_ppwm/u_ex/reg_value_q[0] ),
    .A_N(\u_ppwm/global_counter_high[10] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_497_  (.Y(\u_ppwm/u_ex/_089_ ),
    .B(net383),
    .A_N(\u_ppwm/global_counter_high[13] ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_498_  (.B1(\u_ppwm/u_ex/_089_ ),
    .Y(\u_ppwm/u_ex/_090_ ),
    .A1(\u_ppwm/u_ex/_378_ ),
    .A2(\u_ppwm/global_counter_high[12] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_499_  (.Y(\u_ppwm/u_ex/_091_ ),
    .B(net385),
    .A_N(\u_ppwm/global_counter_high[11] ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_500_  (.A1(\u_ppwm/u_ex/_088_ ),
    .A2(\u_ppwm/u_ex/_091_ ),
    .Y(\u_ppwm/u_ex/_092_ ),
    .B1(\u_ppwm/u_ex/_087_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_501_  (.A(net384),
    .B_N(\u_ppwm/global_counter_high[12] ),
    .Y(\u_ppwm/u_ex/_093_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_502_  (.A(net383),
    .B_N(\u_ppwm/global_counter_high[13] ),
    .Y(\u_ppwm/u_ex/_094_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_503_  (.B2(\u_ppwm/u_ex/_093_ ),
    .C1(\u_ppwm/u_ex/_094_ ),
    .B1(\u_ppwm/u_ex/_089_ ),
    .A1(\u_ppwm/u_ex/_376_ ),
    .Y(\u_ppwm/u_ex/_095_ ),
    .A2(\u_ppwm/global_counter_high[14] ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_504_  (.B1(\u_ppwm/u_ex/_095_ ),
    .Y(\u_ppwm/u_ex/_096_ ),
    .A1(\u_ppwm/u_ex/_090_ ),
    .A2(\u_ppwm/u_ex/_092_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_505_  (.Y(\u_ppwm/u_ex/_097_ ),
    .B1(\u_ppwm/u_ex/_086_ ),
    .B2(\u_ppwm/u_ex/_096_ ),
    .A2(\u_ppwm/global_counter_high[15] ),
    .A1(\u_ppwm/u_ex/_375_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_506_  (.Y(\u_ppwm/u_ex/_098_ ),
    .A(net380),
    .B(\u_ppwm/u_ex/_029_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_507_  (.B1(\u_ppwm/u_ex/_098_ ),
    .Y(\u_ppwm/u_ex/_099_ ),
    .A1(\u_ppwm/u_ex/_375_ ),
    .A2(\u_ppwm/global_counter_high[15] ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_508_  (.B1(\u_ppwm/u_ex/_085_ ),
    .Y(\u_ppwm/u_ex/_100_ ),
    .A1(\u_ppwm/u_ex/_097_ ),
    .A2(\u_ppwm/u_ex/_099_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_509_  (.A(net378),
    .B_N(\u_ppwm/global_counter_high[19] ),
    .Y(\u_ppwm/u_ex/_101_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_510_  (.Y(\u_ppwm/u_ex/_102_ ),
    .B(\u_ppwm/u_ex/reg_value_q[9] ),
    .A_N(\u_ppwm/global_counter_high[19] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_511_  (.Y(\u_ppwm/u_ex/_103_ ),
    .B(\u_ppwm/u_ex/_102_ ),
    .A_N(\u_ppwm/u_ex/_101_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_512_  (.A(\u_ppwm/global_counter_high[18] ),
    .B_N(net379),
    .Y(\u_ppwm/u_ex/_104_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_513_  (.A(\u_ppwm/u_ex/_373_ ),
    .B(\u_ppwm/global_counter_high[17] ),
    .Y(\u_ppwm/u_ex/_105_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_514_  (.A(net379),
    .B_N(\u_ppwm/global_counter_high[18] ),
    .Y(\u_ppwm/u_ex/_106_ ));
 sg13g2_nor4_1 \u_ppwm/u_ex/_515_  (.A(\u_ppwm/u_ex/_103_ ),
    .B(\u_ppwm/u_ex/_104_ ),
    .C(\u_ppwm/u_ex/_105_ ),
    .D(\u_ppwm/u_ex/_106_ ),
    .Y(\u_ppwm/u_ex/_107_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_516_  (.A1(\u_ppwm/u_ex/_102_ ),
    .A2(\u_ppwm/u_ex/_106_ ),
    .Y(\u_ppwm/u_ex/_108_ ),
    .B1(\u_ppwm/u_ex/_101_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_517_  (.B(\u_ppwm/u_ex/_044_ ),
    .C(\u_ppwm/u_ex/_108_ ),
    .A(net324),
    .Y(\u_ppwm/u_ex/_109_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_518_  (.A1(\u_ppwm/u_ex/_100_ ),
    .A2(\u_ppwm/u_ex/_107_ ),
    .Y(\u_ppwm/u_ex/_110_ ),
    .B1(\u_ppwm/u_ex/_109_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_519_  (.Y(\u_ppwm/u_ex/_111_ ),
    .A(\u_ppwm/u_ex/_373_ ),
    .B(net388));
 sg13g2_nor2_1 \u_ppwm/u_ex/_520_  (.A(\u_ppwm/u_ex/_374_ ),
    .B(net389),
    .Y(\u_ppwm/u_ex/_112_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_521_  (.A(net385),
    .B_N(net399),
    .Y(\u_ppwm/u_ex/_113_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_522_  (.Y(\u_ppwm/u_ex/_114_ ),
    .B(\u_ppwm/u_ex/reg_value_q[0] ),
    .A_N(\u_ppwm/pwm_value[0] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_523_  (.Y(\u_ppwm/u_ex/_115_ ),
    .B(net383),
    .A_N(net394));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_524_  (.B1(\u_ppwm/u_ex/_115_ ),
    .Y(\u_ppwm/u_ex/_116_ ),
    .A1(\u_ppwm/u_ex/_378_ ),
    .A2(net396));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_525_  (.Y(\u_ppwm/u_ex/_117_ ),
    .B(net385),
    .A_N(net399));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_526_  (.A1(\u_ppwm/u_ex/_114_ ),
    .A2(\u_ppwm/u_ex/_117_ ),
    .Y(\u_ppwm/u_ex/_118_ ),
    .B1(\u_ppwm/u_ex/_113_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_527_  (.Y(\u_ppwm/u_ex/_119_ ),
    .B1(net397),
    .B2(\u_ppwm/u_ex/_378_ ),
    .A2(net394),
    .A1(\u_ppwm/u_ex/_377_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_528_  (.B1(\u_ppwm/u_ex/_119_ ),
    .Y(\u_ppwm/u_ex/_120_ ),
    .A1(\u_ppwm/u_ex/_116_ ),
    .A2(\u_ppwm/u_ex/_118_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_529_  (.A(net384),
    .B(\u_ppwm/u_ex/_383_ ),
    .C(\u_ppwm/u_ex/_115_ ),
    .Y(\u_ppwm/u_ex/_121_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_530_  (.Y(\u_ppwm/u_ex/_122_ ),
    .B(net393),
    .A_N(net382));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_531_  (.B1(\u_ppwm/u_ex/_122_ ),
    .Y(\u_ppwm/u_ex/_123_ ),
    .A1(net381),
    .A2(\u_ppwm/u_ex/_381_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_532_  (.Y(\u_ppwm/u_ex/_124_ ),
    .B(net381),
    .A_N(net391));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_533_  (.B1(\u_ppwm/u_ex/_124_ ),
    .Y(\u_ppwm/u_ex/_125_ ),
    .A1(\u_ppwm/u_ex/_376_ ),
    .A2(net393));
 sg13g2_nor3_1 \u_ppwm/u_ex/_534_  (.A(\u_ppwm/u_ex/_121_ ),
    .B(\u_ppwm/u_ex/_123_ ),
    .C(\u_ppwm/u_ex/_125_ ),
    .Y(\u_ppwm/u_ex/_126_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_535_  (.A(net380),
    .B_N(net390),
    .Y(\u_ppwm/u_ex/_127_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_536_  (.B2(\u_ppwm/u_ex/_120_ ),
    .C1(\u_ppwm/u_ex/_127_ ),
    .B1(\u_ppwm/u_ex/_126_ ),
    .A1(\u_ppwm/u_ex/_123_ ),
    .Y(\u_ppwm/u_ex/_128_ ),
    .A2(\u_ppwm/u_ex/_124_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_537_  (.B1(\u_ppwm/u_ex/_111_ ),
    .Y(\u_ppwm/u_ex/_129_ ),
    .A1(\u_ppwm/u_ex/_112_ ),
    .A2(\u_ppwm/u_ex/_128_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_538_  (.A(net378),
    .B(\u_ppwm/u_ex/_379_ ),
    .Y(\u_ppwm/u_ex/_130_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_539_  (.Y(\u_ppwm/u_ex/_131_ ),
    .A(net378),
    .B(\u_ppwm/pwm_value[9] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_540_  (.Y(\u_ppwm/u_ex/_132_ ),
    .B(\u_ppwm/u_ex/reg_value_q[7] ),
    .A_N(net387));
 sg13g2_nor2_1 \u_ppwm/u_ex/_541_  (.A(net379),
    .B(\u_ppwm/u_ex/_380_ ),
    .Y(\u_ppwm/u_ex/_133_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_542_  (.Y(\u_ppwm/u_ex/_134_ ),
    .A(net379),
    .B(net386));
 sg13g2_nand4_1 \u_ppwm/u_ex/_543_  (.B(\u_ppwm/u_ex/_131_ ),
    .C(\u_ppwm/u_ex/_132_ ),
    .A(\u_ppwm/u_ex/_129_ ),
    .Y(\u_ppwm/u_ex/_135_ ),
    .D(\u_ppwm/u_ex/_134_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_544_  (.A(net327),
    .B(\u_ppwm/u_ex/_386_ ),
    .C(net324),
    .Y(\u_ppwm/u_ex/_136_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_545_  (.A1(\u_ppwm/u_ex/_131_ ),
    .A2(\u_ppwm/u_ex/_133_ ),
    .Y(\u_ppwm/u_ex/_137_ ),
    .B1(\u_ppwm/u_ex/_130_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_546_  (.A(\u_ppwm/u_ex/_136_ ),
    .B(\u_ppwm/u_ex/_137_ ),
    .X(\u_ppwm/u_ex/_138_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_547_  (.A1(\u_ppwm/u_ex/_135_ ),
    .A2(\u_ppwm/u_ex/_138_ ),
    .Y(\u_ppwm/u_ex/_139_ ),
    .B1(\u_ppwm/u_ex/_110_ ));
 sg13g2_and4_1 \u_ppwm/u_ex/_548_  (.A(net377),
    .B(\u_ppwm/instr[2] ),
    .C(\u_ppwm/u_ex/_385_ ),
    .D(\u_ppwm/instr[1] ),
    .X(\u_ppwm/u_ex/_140_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_549_  (.Y(\u_ppwm/u_ex/_141_ ),
    .B(\u_ppwm/global_counter_high[1] ),
    .A_N(net398));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_550_  (.A(\u_ppwm/global_counter_high[0] ),
    .B_N(\u_ppwm/pwm_value[0] ),
    .Y(\u_ppwm/u_ex/_142_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_551_  (.A(\u_ppwm/global_counter_high[1] ),
    .B_N(net398),
    .Y(\u_ppwm/u_ex/_143_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_552_  (.B2(\u_ppwm/u_ex/_142_ ),
    .C1(\u_ppwm/u_ex/_143_ ),
    .B1(\u_ppwm/u_ex/_141_ ),
    .A1(net397),
    .Y(\u_ppwm/u_ex/_144_ ),
    .A2(\u_ppwm/u_ex/_039_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_553_  (.Y(\u_ppwm/u_ex/_145_ ),
    .B(\u_ppwm/global_counter_high[3] ),
    .A_N(net395));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_554_  (.B1(\u_ppwm/u_ex/_145_ ),
    .Y(\u_ppwm/u_ex/_146_ ),
    .A1(net397),
    .A2(\u_ppwm/u_ex/_039_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_555_  (.A(\u_ppwm/global_counter_high[5] ),
    .B_N(\u_ppwm/pwm_value[5] ),
    .Y(\u_ppwm/u_ex/_147_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_556_  (.A(\u_ppwm/global_counter_high[3] ),
    .B_N(net395),
    .Y(\u_ppwm/u_ex/_148_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_557_  (.B(\u_ppwm/global_counter_high[4] ),
    .A(net393),
    .X(\u_ppwm/u_ex/_149_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_558_  (.A(\u_ppwm/u_ex/_147_ ),
    .B(\u_ppwm/u_ex/_148_ ),
    .C(\u_ppwm/u_ex/_149_ ),
    .Y(\u_ppwm/u_ex/_150_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_559_  (.B1(\u_ppwm/u_ex/_150_ ),
    .Y(\u_ppwm/u_ex/_151_ ),
    .A1(\u_ppwm/u_ex/_144_ ),
    .A2(\u_ppwm/u_ex/_146_ ));
 sg13g2_nor3_1 \u_ppwm/u_ex/_560_  (.A(net393),
    .B(\u_ppwm/u_ex/_037_ ),
    .C(\u_ppwm/u_ex/_147_ ),
    .Y(\u_ppwm/u_ex/_152_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_561_  (.A1(\u_ppwm/u_ex/_381_ ),
    .A2(\u_ppwm/global_counter_high[5] ),
    .Y(\u_ppwm/u_ex/_153_ ),
    .B1(\u_ppwm/u_ex/_152_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_562_  (.A(net390),
    .B(\u_ppwm/u_ex/_036_ ),
    .Y(\u_ppwm/u_ex/_154_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_563_  (.Y(\u_ppwm/u_ex/_155_ ),
    .A(net387),
    .B(\u_ppwm/u_ex/_035_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_564_  (.B1(\u_ppwm/u_ex/_155_ ),
    .Y(\u_ppwm/u_ex/_156_ ),
    .A1(net390),
    .A2(\u_ppwm/u_ex/_036_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_565_  (.B2(\u_ppwm/u_ex/_153_ ),
    .C1(\u_ppwm/u_ex/_156_ ),
    .B1(\u_ppwm/u_ex/_151_ ),
    .A1(net390),
    .Y(\u_ppwm/u_ex/_157_ ),
    .A2(\u_ppwm/u_ex/_036_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_566_  (.A(net388),
    .B(\u_ppwm/u_ex/_035_ ),
    .Y(\u_ppwm/u_ex/_158_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_567_  (.B1(\u_ppwm/u_ex/_155_ ),
    .Y(\u_ppwm/u_ex/_159_ ),
    .A1(\u_ppwm/u_ex/_154_ ),
    .A2(\u_ppwm/u_ex/_158_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_568_  (.B1(\u_ppwm/u_ex/_159_ ),
    .Y(\u_ppwm/u_ex/_160_ ),
    .A1(\u_ppwm/pwm_value[8] ),
    .A2(\u_ppwm/u_ex/_034_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_569_  (.Y(\u_ppwm/u_ex/_161_ ),
    .B1(\u_ppwm/u_ex/_034_ ),
    .B2(\u_ppwm/pwm_value[8] ),
    .A2(\u_ppwm/u_ex/_033_ ),
    .A1(\u_ppwm/pwm_value[9] ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_570_  (.B1(\u_ppwm/u_ex/_161_ ),
    .Y(\u_ppwm/u_ex/_162_ ),
    .A1(\u_ppwm/u_ex/_157_ ),
    .A2(\u_ppwm/u_ex/_160_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_571_  (.A(net327),
    .B(net325),
    .Y(\u_ppwm/u_ex/_163_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_572_  (.A1(\u_ppwm/u_ex/_379_ ),
    .A2(\u_ppwm/global_counter_high[9] ),
    .Y(\u_ppwm/u_ex/_164_ ),
    .B1(net324));
 sg13g2_nand3_1 \u_ppwm/u_ex/_573_  (.B(\u_ppwm/u_ex/_163_ ),
    .C(\u_ppwm/u_ex/_164_ ),
    .A(\u_ppwm/u_ex/_162_ ),
    .Y(\u_ppwm/u_ex/_165_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_574_  (.Y(\u_ppwm/u_ex/_166_ ),
    .B1(\u_ppwm/global_counter_high[14] ),
    .B2(\u_ppwm/u_ex/_382_ ),
    .A2(\u_ppwm/global_counter_high[15] ),
    .A1(\u_ppwm/u_ex/_381_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_575_  (.Y(\u_ppwm/u_ex/_167_ ),
    .B(\u_ppwm/global_counter_high[11] ),
    .A_N(net399));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_576_  (.A(\u_ppwm/global_counter_high[10] ),
    .B_N(\u_ppwm/pwm_value[0] ),
    .Y(\u_ppwm/u_ex/_168_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_577_  (.A(\u_ppwm/global_counter_high[11] ),
    .B_N(net399),
    .Y(\u_ppwm/u_ex/_169_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_578_  (.B2(\u_ppwm/u_ex/_168_ ),
    .C1(\u_ppwm/u_ex/_169_ ),
    .B1(\u_ppwm/u_ex/_167_ ),
    .A1(net397),
    .Y(\u_ppwm/u_ex/_170_ ),
    .A2(\u_ppwm/u_ex/_032_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_579_  (.Y(\u_ppwm/u_ex/_171_ ),
    .B(\u_ppwm/global_counter_high[13] ),
    .A_N(net395));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_580_  (.B1(\u_ppwm/u_ex/_171_ ),
    .Y(\u_ppwm/u_ex/_172_ ),
    .A1(net397),
    .A2(\u_ppwm/u_ex/_032_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_581_  (.Y(\u_ppwm/u_ex/_173_ ),
    .B1(\u_ppwm/u_ex/_031_ ),
    .B2(net395),
    .A2(\u_ppwm/u_ex/_030_ ),
    .A1(net393));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_582_  (.B1(\u_ppwm/u_ex/_173_ ),
    .Y(\u_ppwm/u_ex/_174_ ),
    .A1(\u_ppwm/u_ex/_170_ ),
    .A2(\u_ppwm/u_ex/_172_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_583_  (.A(\u_ppwm/u_ex/_381_ ),
    .B(\u_ppwm/global_counter_high[15] ),
    .Y(\u_ppwm/u_ex/_175_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_584_  (.B2(\u_ppwm/u_ex/_174_ ),
    .C1(\u_ppwm/u_ex/_175_ ),
    .B1(\u_ppwm/u_ex/_166_ ),
    .A1(net390),
    .Y(\u_ppwm/u_ex/_176_ ),
    .A2(\u_ppwm/u_ex/_029_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_585_  (.Y(\u_ppwm/u_ex/_177_ ),
    .B(\u_ppwm/global_counter_high[17] ),
    .A_N(net388));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_586_  (.B1(\u_ppwm/u_ex/_177_ ),
    .Y(\u_ppwm/u_ex/_178_ ),
    .A1(net390),
    .A2(\u_ppwm/u_ex/_029_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_587_  (.Y(\u_ppwm/u_ex/_179_ ),
    .B1(\u_ppwm/global_counter_high[18] ),
    .B2(\u_ppwm/u_ex/_380_ ),
    .A2(\u_ppwm/global_counter_high[19] ),
    .A1(\u_ppwm/u_ex/_379_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_588_  (.Y(\u_ppwm/u_ex/_180_ ),
    .B(\u_ppwm/pwm_value[9] ),
    .A_N(\u_ppwm/global_counter_high[19] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_589_  (.Y(\u_ppwm/u_ex/_181_ ),
    .B(net388),
    .A_N(\u_ppwm/global_counter_high[17] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_590_  (.Y(\u_ppwm/u_ex/_182_ ),
    .B(\u_ppwm/pwm_value[8] ),
    .A_N(\u_ppwm/global_counter_high[18] ));
 sg13g2_and4_1 \u_ppwm/u_ex/_591_  (.A(\u_ppwm/u_ex/_179_ ),
    .B(\u_ppwm/u_ex/_180_ ),
    .C(\u_ppwm/u_ex/_181_ ),
    .D(\u_ppwm/u_ex/_182_ ),
    .X(\u_ppwm/u_ex/_183_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_592_  (.B1(\u_ppwm/u_ex/_183_ ),
    .Y(\u_ppwm/u_ex/_184_ ),
    .A1(\u_ppwm/u_ex/_176_ ),
    .A2(\u_ppwm/u_ex/_178_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_593_  (.Y(\u_ppwm/u_ex/_185_ ),
    .B(\u_ppwm/u_ex/_180_ ),
    .A_N(\u_ppwm/u_ex/_179_ ));
 sg13g2_nand4_1 \u_ppwm/u_ex/_594_  (.B(\u_ppwm/u_ex/_163_ ),
    .C(\u_ppwm/u_ex/_184_ ),
    .A(net324),
    .Y(\u_ppwm/u_ex/_186_ ),
    .D(\u_ppwm/u_ex/_185_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_595_  (.A(net380),
    .B(\u_ppwm/u_ex/_036_ ),
    .Y(\u_ppwm/u_ex/_187_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_596_  (.Y(\u_ppwm/u_ex/_188_ ),
    .B(\u_ppwm/global_counter_high[1] ),
    .A_N(net385));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_597_  (.A(\u_ppwm/global_counter_high[0] ),
    .B_N(\u_ppwm/u_ex/reg_value_q[0] ),
    .Y(\u_ppwm/u_ex/_189_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_598_  (.A(\u_ppwm/global_counter_high[1] ),
    .B_N(net385),
    .Y(\u_ppwm/u_ex/_190_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_599_  (.B2(\u_ppwm/u_ex/_189_ ),
    .C1(\u_ppwm/u_ex/_190_ ),
    .B1(\u_ppwm/u_ex/_188_ ),
    .A1(net384),
    .Y(\u_ppwm/u_ex/_191_ ),
    .A2(\u_ppwm/u_ex/_039_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_600_  (.B2(\u_ppwm/u_ex/_378_ ),
    .C1(\u_ppwm/u_ex/_191_ ),
    .B1(\u_ppwm/global_counter_high[2] ),
    .A1(\u_ppwm/u_ex/_377_ ),
    .Y(\u_ppwm/u_ex/_192_ ),
    .A2(\u_ppwm/global_counter_high[3] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_601_  (.Y(\u_ppwm/u_ex/_193_ ),
    .B(net381),
    .A_N(\u_ppwm/global_counter_high[5] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_602_  (.Y(\u_ppwm/u_ex/_194_ ),
    .B(\u_ppwm/global_counter_high[4] ),
    .A_N(net382));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_603_  (.Y(\u_ppwm/u_ex/_195_ ),
    .B1(\u_ppwm/u_ex/_038_ ),
    .B2(net383),
    .A2(\u_ppwm/u_ex/_037_ ),
    .A1(net382));
 sg13g2_nand3_1 \u_ppwm/u_ex/_604_  (.B(\u_ppwm/u_ex/_194_ ),
    .C(\u_ppwm/u_ex/_195_ ),
    .A(\u_ppwm/u_ex/_193_ ),
    .Y(\u_ppwm/u_ex/_196_ ));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_605_  (.A(\u_ppwm/u_ex/_194_ ),
    .B_N(\u_ppwm/u_ex/_193_ ),
    .Y(\u_ppwm/u_ex/_197_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_606_  (.A1(\u_ppwm/u_ex/_375_ ),
    .A2(\u_ppwm/global_counter_high[5] ),
    .Y(\u_ppwm/u_ex/_198_ ),
    .B1(\u_ppwm/u_ex/_197_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_607_  (.B1(\u_ppwm/u_ex/_198_ ),
    .Y(\u_ppwm/u_ex/_199_ ),
    .A1(\u_ppwm/u_ex/_192_ ),
    .A2(\u_ppwm/u_ex/_196_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_608_  (.Y(\u_ppwm/u_ex/_200_ ),
    .A(net380),
    .B(\u_ppwm/u_ex/_036_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_609_  (.B2(\u_ppwm/u_ex/_200_ ),
    .C1(\u_ppwm/u_ex/_187_ ),
    .B1(\u_ppwm/u_ex/_199_ ),
    .A1(\u_ppwm/u_ex/_373_ ),
    .Y(\u_ppwm/u_ex/_201_ ),
    .A2(\u_ppwm/global_counter_high[7] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_610_  (.Y(\u_ppwm/u_ex/_202_ ),
    .B(\u_ppwm/global_counter_high[9] ),
    .A_N(net378));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_611_  (.B1(\u_ppwm/u_ex/_202_ ),
    .Y(\u_ppwm/u_ex/_203_ ),
    .A1(net379),
    .A2(\u_ppwm/u_ex/_034_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_612_  (.Y(\u_ppwm/u_ex/_204_ ),
    .A(net378),
    .B(\u_ppwm/u_ex/_033_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_613_  (.Y(\u_ppwm/u_ex/_205_ ),
    .B1(\u_ppwm/u_ex/_035_ ),
    .B2(\u_ppwm/u_ex/reg_value_q[7] ),
    .A2(\u_ppwm/u_ex/_034_ ),
    .A1(net379));
 sg13g2_nand3b_1 \u_ppwm/u_ex/_614_  (.B(\u_ppwm/u_ex/_204_ ),
    .C(\u_ppwm/u_ex/_205_ ),
    .Y(\u_ppwm/u_ex/_206_ ),
    .A_N(\u_ppwm/u_ex/_203_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_615_  (.A1(\u_ppwm/u_ex/_203_ ),
    .A2(\u_ppwm/u_ex/_204_ ),
    .Y(\u_ppwm/u_ex/_207_ ),
    .B1(\u_ppwm/u_ex/_045_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_616_  (.B1(\u_ppwm/u_ex/_207_ ),
    .Y(\u_ppwm/u_ex/_208_ ),
    .A1(\u_ppwm/u_ex/_201_ ),
    .A2(\u_ppwm/u_ex/_206_ ));
 sg13g2_and4_1 \u_ppwm/u_ex/_617_  (.A(\u_ppwm/u_ex/_140_ ),
    .B(\u_ppwm/u_ex/_165_ ),
    .C(\u_ppwm/u_ex/_186_ ),
    .D(\u_ppwm/u_ex/_208_ ),
    .X(\u_ppwm/u_ex/_209_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_618_  (.B1(net439),
    .Y(\u_ppwm/u_ex/_210_ ),
    .A1(net627),
    .A2(\u_ppwm/u_ex/_140_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_619_  (.A1(\u_ppwm/u_ex/_139_ ),
    .A2(\u_ppwm/u_ex/_209_ ),
    .Y(\u_ppwm/u_ex/_007_ ),
    .B1(net628));
 sg13g2_nand2_1 \u_ppwm/u_ex/_620_  (.Y(\u_ppwm/u_ex/_211_ ),
    .A(net377),
    .B(\u_ppwm/u_ex/_046_ ));
 sg13g2_nor2_2 \u_ppwm/u_ex/_621_  (.A(\u_ppwm/instr[2] ),
    .B(\u_ppwm/u_ex/_211_ ),
    .Y(\u_ppwm/u_ex/_212_ ));
 sg13g2_nor3_2 \u_ppwm/u_ex/_622_  (.A(\u_ppwm/instr[2] ),
    .B(net327),
    .C(\u_ppwm/u_ex/_211_ ),
    .Y(\u_ppwm/u_ex/_213_ ));
 sg13g2_nand2b_2 \u_ppwm/u_ex/_623_  (.Y(\u_ppwm/u_ex/_214_ ),
    .B(\u_ppwm/u_ex/_212_ ),
    .A_N(net327));
 sg13g2_nand2b_2 \u_ppwm/u_ex/_624_  (.Y(\u_ppwm/u_ex/_215_ ),
    .B(\u_ppwm/instr[1] ),
    .A_N(\u_ppwm/instr[2] ));
 sg13g2_nor2_2 \u_ppwm/u_ex/_625_  (.A(\u_ppwm/instr[0] ),
    .B(net317),
    .Y(\u_ppwm/u_ex/_216_ ));
 sg13g2_nand2b_2 \u_ppwm/u_ex/_626_  (.Y(\u_ppwm/u_ex/_217_ ),
    .B(\u_ppwm/u_ex/_385_ ),
    .A_N(net317));
 sg13g2_and2_1 \u_ppwm/u_ex/_627_  (.A(\u_ppwm/pwm_value[0] ),
    .B(net325),
    .X(\u_ppwm/u_ex/_218_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_628_  (.B1(net310),
    .Y(\u_ppwm/u_ex/_219_ ),
    .A1(net315),
    .A2(\u_ppwm/u_ex/_218_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_629_  (.B1(\u_ppwm/u_ex/_219_ ),
    .Y(\u_ppwm/u_ex/_220_ ),
    .A1(net649),
    .A2(net325));
 sg13g2_nor3_2 \u_ppwm/u_ex/_630_  (.A(\u_ppwm/u_ex/_385_ ),
    .B(net325),
    .C(net317),
    .Y(\u_ppwm/u_ex/_221_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_631_  (.Y(\u_ppwm/u_ex/_222_ ),
    .B1(net314),
    .B2(net398),
    .A2(net317),
    .A1(net325));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_632_  (.B1(net439),
    .Y(\u_ppwm/u_ex/_223_ ),
    .A1(net649),
    .A2(\u_ppwm/u_ex/_213_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_633_  (.A1(\u_ppwm/u_ex/_220_ ),
    .A2(\u_ppwm/u_ex/_222_ ),
    .Y(\u_ppwm/u_ex/_008_ ),
    .B1(\u_ppwm/u_ex/_223_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_634_  (.A(net398),
    .B(net323),
    .X(\u_ppwm/u_ex/_224_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_635_  (.B(net323),
    .A(net398),
    .X(\u_ppwm/u_ex/_225_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_636_  (.B(\u_ppwm/u_ex/_225_ ),
    .A(\u_ppwm/u_ex/_218_ ),
    .X(\u_ppwm/u_ex/_226_ ));
 sg13g2_nor3_2 \u_ppwm/u_ex/_637_  (.A(\u_ppwm/u_ex/_385_ ),
    .B(\u_ppwm/u_ex/_386_ ),
    .C(net317),
    .Y(\u_ppwm/u_ex/_227_ ));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_638_  (.Y(\u_ppwm/u_ex/_228_ ),
    .B1(net316),
    .B2(\u_ppwm/u_ex/_226_ ),
    .A2(net317),
    .A1(net323));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_639_  (.B2(net649),
    .C1(net309),
    .B1(net311),
    .A1(net396),
    .Y(\u_ppwm/u_ex/_229_ ),
    .A2(net313));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_640_  (.B1(net426),
    .Y(\u_ppwm/u_ex/_230_ ),
    .A1(net398),
    .A2(\u_ppwm/u_ex/_213_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_641_  (.A1(\u_ppwm/u_ex/_228_ ),
    .A2(\u_ppwm/u_ex/_229_ ),
    .Y(\u_ppwm/u_ex/_009_ ),
    .B1(\u_ppwm/u_ex/_230_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_642_  (.A1(\u_ppwm/u_ex/_218_ ),
    .A2(\u_ppwm/u_ex/_225_ ),
    .Y(\u_ppwm/u_ex/_231_ ),
    .B1(\u_ppwm/u_ex/_224_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_643_  (.Y(\u_ppwm/u_ex/_232_ ),
    .A(net396),
    .B(net319));
 sg13g2_nor2_1 \u_ppwm/u_ex/_644_  (.A(\u_ppwm/u_ex/_231_ ),
    .B(\u_ppwm/u_ex/_232_ ),
    .Y(\u_ppwm/u_ex/_233_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_645_  (.A1(\u_ppwm/u_ex/_231_ ),
    .A2(\u_ppwm/u_ex/_232_ ),
    .Y(\u_ppwm/u_ex/_234_ ),
    .B1(net315));
 sg13g2_nor2b_1 \u_ppwm/u_ex/_646_  (.A(\u_ppwm/u_ex/_233_ ),
    .B_N(\u_ppwm/u_ex/_234_ ),
    .Y(\u_ppwm/u_ex/_235_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_647_  (.Y(\u_ppwm/u_ex/_236_ ),
    .A(net320),
    .B(net317));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_648_  (.Y(\u_ppwm/u_ex/_237_ ),
    .B1(net312),
    .B2(net398),
    .A2(net314),
    .A1(net394));
 sg13g2_nand3_1 \u_ppwm/u_ex/_649_  (.B(\u_ppwm/u_ex/_236_ ),
    .C(\u_ppwm/u_ex/_237_ ),
    .A(net310),
    .Y(\u_ppwm/u_ex/_238_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_650_  (.B1(net439),
    .Y(\u_ppwm/u_ex/_239_ ),
    .A1(\u_ppwm/u_ex/_235_ ),
    .A2(\u_ppwm/u_ex/_238_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_651_  (.A1(\u_ppwm/u_ex/_383_ ),
    .A2(net309),
    .Y(\u_ppwm/u_ex/_010_ ),
    .B1(\u_ppwm/u_ex/_239_ ));
 sg13g2_xor2_1 \u_ppwm/u_ex/_652_  (.B(net319),
    .A(net394),
    .X(\u_ppwm/u_ex/_240_ ));
 sg13g2_a21o_1 \u_ppwm/u_ex/_653_  (.A2(net320),
    .A1(net396),
    .B1(\u_ppwm/u_ex/_233_ ),
    .X(\u_ppwm/u_ex/_241_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_654_  (.A1(\u_ppwm/u_ex/_240_ ),
    .A2(\u_ppwm/u_ex/_241_ ),
    .Y(\u_ppwm/u_ex/_242_ ),
    .B1(net315));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_655_  (.B1(\u_ppwm/u_ex/_242_ ),
    .Y(\u_ppwm/u_ex/_243_ ),
    .A1(\u_ppwm/u_ex/_240_ ),
    .A2(\u_ppwm/u_ex/_241_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_656_  (.B2(net396),
    .C1(\u_ppwm/u_ex/_214_ ),
    .B1(net311),
    .A1(net392),
    .Y(\u_ppwm/u_ex/_244_ ),
    .A2(net313));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_657_  (.B1(net427),
    .Y(\u_ppwm/u_ex/_245_ ),
    .A1(net394),
    .A2(\u_ppwm/u_ex/_213_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_658_  (.A1(\u_ppwm/u_ex/_243_ ),
    .A2(\u_ppwm/u_ex/_244_ ),
    .Y(\u_ppwm/u_ex/_011_ ),
    .B1(\u_ppwm/u_ex/_245_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_659_  (.Y(\u_ppwm/u_ex/_246_ ),
    .B(\u_ppwm/u_ex/_240_ ),
    .A_N(\u_ppwm/u_ex/_232_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_660_  (.B1(net319),
    .Y(\u_ppwm/u_ex/_247_ ),
    .A1(net394),
    .A2(net396));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_661_  (.B1(\u_ppwm/u_ex/_247_ ),
    .Y(\u_ppwm/u_ex/_248_ ),
    .A1(\u_ppwm/u_ex/_231_ ),
    .A2(\u_ppwm/u_ex/_246_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_662_  (.Y(\u_ppwm/u_ex/_249_ ),
    .A(net392),
    .B(net318));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_663_  (.Y(\u_ppwm/u_ex/_250_ ),
    .A(net392),
    .B(net318));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_664_  (.Y(\u_ppwm/u_ex/_251_ ),
    .B(\u_ppwm/u_ex/_248_ ),
    .A_N(\u_ppwm/u_ex/_250_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_665_  (.Y(\u_ppwm/u_ex/_252_ ),
    .B(\u_ppwm/u_ex/_250_ ),
    .A_N(\u_ppwm/u_ex/_248_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_666_  (.B(\u_ppwm/u_ex/_251_ ),
    .C(\u_ppwm/u_ex/_252_ ),
    .A(net316),
    .Y(\u_ppwm/u_ex/_253_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_667_  (.B2(net394),
    .C1(net309),
    .B1(net311),
    .A1(net391),
    .Y(\u_ppwm/u_ex/_254_ ),
    .A2(net313));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_668_  (.B1(net425),
    .Y(\u_ppwm/u_ex/_255_ ),
    .A1(net392),
    .A2(net310));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_669_  (.A1(\u_ppwm/u_ex/_253_ ),
    .A2(\u_ppwm/u_ex/_254_ ),
    .Y(\u_ppwm/u_ex/_012_ ),
    .B1(\u_ppwm/u_ex/_255_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_670_  (.Y(\u_ppwm/u_ex/_256_ ),
    .A(net391),
    .B(net318));
 sg13g2_nand3_1 \u_ppwm/u_ex/_671_  (.B(\u_ppwm/u_ex/_251_ ),
    .C(\u_ppwm/u_ex/_256_ ),
    .A(\u_ppwm/u_ex/_249_ ),
    .Y(\u_ppwm/u_ex/_257_ ));
 sg13g2_a21o_1 \u_ppwm/u_ex/_672_  (.A2(\u_ppwm/u_ex/_251_ ),
    .A1(\u_ppwm/u_ex/_249_ ),
    .B1(\u_ppwm/u_ex/_256_ ),
    .X(\u_ppwm/u_ex/_258_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_673_  (.B(\u_ppwm/u_ex/_257_ ),
    .C(\u_ppwm/u_ex/_258_ ),
    .A(net316),
    .Y(\u_ppwm/u_ex/_259_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_674_  (.B2(net392),
    .C1(net309),
    .B1(net311),
    .A1(net389),
    .Y(\u_ppwm/u_ex/_260_ ),
    .A2(net313));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_675_  (.B1(net425),
    .Y(\u_ppwm/u_ex/_261_ ),
    .A1(net391),
    .A2(net310));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_676_  (.A1(\u_ppwm/u_ex/_259_ ),
    .A2(\u_ppwm/u_ex/_260_ ),
    .Y(\u_ppwm/u_ex/_013_ ),
    .B1(\u_ppwm/u_ex/_261_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_677_  (.Y(\u_ppwm/u_ex/_262_ ),
    .A(net389),
    .B(net318));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_678_  (.Y(\u_ppwm/u_ex/_263_ ),
    .A(net389),
    .B(net318));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_679_  (.B1(net318),
    .Y(\u_ppwm/u_ex/_264_ ),
    .A1(net391),
    .A2(net392));
 sg13g2_inv_1 \u_ppwm/u_ex/_680_  (.Y(\u_ppwm/u_ex/_265_ ),
    .A(\u_ppwm/u_ex/_264_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_681_  (.A(\u_ppwm/u_ex/_250_ ),
    .B(\u_ppwm/u_ex/_256_ ),
    .Y(\u_ppwm/u_ex/_266_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_682_  (.A1(\u_ppwm/u_ex/_248_ ),
    .A2(\u_ppwm/u_ex/_266_ ),
    .Y(\u_ppwm/u_ex/_267_ ),
    .B1(\u_ppwm/u_ex/_265_ ));
 sg13g2_or2_1 \u_ppwm/u_ex/_683_  (.X(\u_ppwm/u_ex/_268_ ),
    .B(\u_ppwm/u_ex/_267_ ),
    .A(\u_ppwm/u_ex/_263_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_684_  (.A1(\u_ppwm/u_ex/_263_ ),
    .A2(\u_ppwm/u_ex/_267_ ),
    .Y(\u_ppwm/u_ex/_269_ ),
    .B1(net315));
 sg13g2_nand2_1 \u_ppwm/u_ex/_685_  (.Y(\u_ppwm/u_ex/_270_ ),
    .A(\u_ppwm/u_ex/_268_ ),
    .B(\u_ppwm/u_ex/_269_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_686_  (.B2(net391),
    .C1(net309),
    .B1(net311),
    .A1(net387),
    .Y(\u_ppwm/u_ex/_271_ ),
    .A2(net313));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_687_  (.B1(net426),
    .Y(\u_ppwm/u_ex/_272_ ),
    .A1(net389),
    .A2(net310));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_688_  (.A1(\u_ppwm/u_ex/_270_ ),
    .A2(\u_ppwm/u_ex/_271_ ),
    .Y(\u_ppwm/u_ex/_014_ ),
    .B1(\u_ppwm/u_ex/_272_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_689_  (.Y(\u_ppwm/u_ex/_273_ ),
    .A(net387),
    .B(net318));
 sg13g2_nand3_1 \u_ppwm/u_ex/_690_  (.B(\u_ppwm/u_ex/_268_ ),
    .C(\u_ppwm/u_ex/_273_ ),
    .A(\u_ppwm/u_ex/_262_ ),
    .Y(\u_ppwm/u_ex/_274_ ));
 sg13g2_a21o_1 \u_ppwm/u_ex/_691_  (.A2(\u_ppwm/u_ex/_268_ ),
    .A1(\u_ppwm/u_ex/_262_ ),
    .B1(\u_ppwm/u_ex/_273_ ),
    .X(\u_ppwm/u_ex/_275_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_692_  (.B(\u_ppwm/u_ex/_274_ ),
    .C(\u_ppwm/u_ex/_275_ ),
    .A(net316),
    .Y(\u_ppwm/u_ex/_276_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_693_  (.B2(net389),
    .C1(net309),
    .B1(net311),
    .A1(net386),
    .Y(\u_ppwm/u_ex/_277_ ),
    .A2(net313));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_694_  (.B1(net426),
    .Y(\u_ppwm/u_ex/_278_ ),
    .A1(net387),
    .A2(net310));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_695_  (.A1(\u_ppwm/u_ex/_276_ ),
    .A2(\u_ppwm/u_ex/_277_ ),
    .Y(\u_ppwm/u_ex/_015_ ),
    .B1(\u_ppwm/u_ex/_278_ ));
 sg13g2_nor4_1 \u_ppwm/u_ex/_696_  (.A(\u_ppwm/u_ex/_250_ ),
    .B(\u_ppwm/u_ex/_256_ ),
    .C(\u_ppwm/u_ex/_263_ ),
    .D(\u_ppwm/u_ex/_273_ ),
    .Y(\u_ppwm/u_ex/_279_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_697_  (.B1(net318),
    .Y(\u_ppwm/u_ex/_280_ ),
    .A1(net387),
    .A2(net389));
 sg13g2_nand2_1 \u_ppwm/u_ex/_698_  (.Y(\u_ppwm/u_ex/_281_ ),
    .A(\u_ppwm/u_ex/_264_ ),
    .B(\u_ppwm/u_ex/_280_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_699_  (.A1(\u_ppwm/u_ex/_248_ ),
    .A2(\u_ppwm/u_ex/_279_ ),
    .Y(\u_ppwm/u_ex/_282_ ),
    .B1(\u_ppwm/u_ex/_281_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_700_  (.Y(\u_ppwm/u_ex/_283_ ),
    .A(net386),
    .B(net319));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_701_  (.Y(\u_ppwm/u_ex/_284_ ),
    .A(net386),
    .B(net319));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_702_  (.A1(\u_ppwm/u_ex/_282_ ),
    .A2(\u_ppwm/u_ex/_284_ ),
    .Y(\u_ppwm/u_ex/_285_ ),
    .B1(net315));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_703_  (.B1(\u_ppwm/u_ex/_285_ ),
    .Y(\u_ppwm/u_ex/_286_ ),
    .A1(\u_ppwm/u_ex/_282_ ),
    .A2(\u_ppwm/u_ex/_284_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_704_  (.B2(net387),
    .C1(net309),
    .B1(net311),
    .A1(net651),
    .Y(\u_ppwm/u_ex/_287_ ),
    .A2(net313));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_705_  (.B1(net426),
    .Y(\u_ppwm/u_ex/_288_ ),
    .A1(net386),
    .A2(net310));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_706_  (.A1(\u_ppwm/u_ex/_286_ ),
    .A2(\u_ppwm/u_ex/_287_ ),
    .Y(\u_ppwm/u_ex/_016_ ),
    .B1(\u_ppwm/u_ex/_288_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_707_  (.B1(\u_ppwm/u_ex/_283_ ),
    .Y(\u_ppwm/u_ex/_289_ ),
    .A1(\u_ppwm/u_ex/_282_ ),
    .A2(\u_ppwm/u_ex/_284_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_708_  (.Y(\u_ppwm/u_ex/_290_ ),
    .A(\u_ppwm/pwm_value[9] ),
    .B(net319));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_709_  (.Y(\u_ppwm/u_ex/_291_ ),
    .A(\u_ppwm/u_ex/_289_ ),
    .B(\u_ppwm/u_ex/_290_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_710_  (.B2(net316),
    .C1(net309),
    .B1(\u_ppwm/u_ex/_291_ ),
    .A1(net386),
    .Y(\u_ppwm/u_ex/_292_ ),
    .A2(net311));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_711_  (.B1(net426),
    .Y(\u_ppwm/u_ex/_293_ ),
    .A1(net651),
    .A2(net310));
 sg13g2_nor2_1 \u_ppwm/u_ex/_712_  (.A(\u_ppwm/u_ex/_292_ ),
    .B(\u_ppwm/u_ex/_293_ ),
    .Y(\u_ppwm/u_ex/_017_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_713_  (.A(net327),
    .B(\u_ppwm/u_ex/_212_ ),
    .X(\u_ppwm/u_ex/_294_ ));
 sg13g2_nand2_2 \u_ppwm/u_ex/_714_  (.Y(\u_ppwm/u_ex/_295_ ),
    .A(net327),
    .B(\u_ppwm/u_ex/_212_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_715_  (.A(\u_ppwm/u_ex/reg_value_q[0] ),
    .B(net325),
    .X(\u_ppwm/u_ex/_296_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_716_  (.Y(\u_ppwm/u_ex/_297_ ),
    .A(net641),
    .B(net326));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_717_  (.B1(net307),
    .Y(\u_ppwm/u_ex/_298_ ),
    .A1(net315),
    .A2(\u_ppwm/u_ex/_296_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_718_  (.B1(\u_ppwm/u_ex/_298_ ),
    .Y(\u_ppwm/u_ex/_299_ ),
    .A1(\u_ppwm/u_ex/reg_value_q[0] ),
    .A2(net326));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_719_  (.Y(\u_ppwm/u_ex/_300_ ),
    .B1(net313),
    .B2(net634),
    .A2(net317),
    .A1(net326));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_720_  (.B1(net442),
    .Y(\u_ppwm/u_ex/_301_ ),
    .A1(\u_ppwm/u_ex/reg_value_q[0] ),
    .A2(net307));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_721_  (.A1(\u_ppwm/u_ex/_299_ ),
    .A2(\u_ppwm/u_ex/_300_ ),
    .Y(\u_ppwm/u_ex/_018_ ),
    .B1(\u_ppwm/u_ex/_301_ ));
 sg13g2_and2_1 \u_ppwm/u_ex/_722_  (.A(net385),
    .B(net323),
    .X(\u_ppwm/u_ex/_302_ ));
 sg13g2_or2_1 \u_ppwm/u_ex/_723_  (.X(\u_ppwm/u_ex/_303_ ),
    .B(net323),
    .A(\u_ppwm/u_ex/reg_value_q[1] ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_724_  (.Y(\u_ppwm/u_ex/_304_ ),
    .B(\u_ppwm/u_ex/_303_ ),
    .A_N(\u_ppwm/u_ex/_302_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_725_  (.B1(net316),
    .Y(\u_ppwm/u_ex/_305_ ),
    .A1(\u_ppwm/u_ex/_297_ ),
    .A2(\u_ppwm/u_ex/_304_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_726_  (.A1(\u_ppwm/u_ex/_297_ ),
    .A2(\u_ppwm/u_ex/_304_ ),
    .Y(\u_ppwm/u_ex/_306_ ),
    .B1(\u_ppwm/u_ex/_305_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_727_  (.A1(net384),
    .A2(net314),
    .Y(\u_ppwm/u_ex/_307_ ),
    .B1(\u_ppwm/u_ex/_295_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_728_  (.B2(net641),
    .C1(\u_ppwm/u_ex/_306_ ),
    .B1(net312),
    .A1(net323),
    .Y(\u_ppwm/u_ex/_308_ ),
    .A2(\u_ppwm/u_ex/_215_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_729_  (.B1(net442),
    .Y(\u_ppwm/u_ex/_309_ ),
    .A1(net634),
    .A2(net307));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_730_  (.A1(\u_ppwm/u_ex/_307_ ),
    .A2(\u_ppwm/u_ex/_308_ ),
    .Y(\u_ppwm/u_ex/_019_ ),
    .B1(\u_ppwm/u_ex/_309_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_731_  (.A1(\u_ppwm/u_ex/_296_ ),
    .A2(\u_ppwm/u_ex/_303_ ),
    .Y(\u_ppwm/u_ex/_310_ ),
    .B1(\u_ppwm/u_ex/_302_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_732_  (.Y(\u_ppwm/u_ex/_311_ ),
    .A(net384),
    .B(net322));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_733_  (.Y(\u_ppwm/u_ex/_312_ ),
    .A(net384),
    .B(net322));
 sg13g2_or2_1 \u_ppwm/u_ex/_734_  (.X(\u_ppwm/u_ex/_313_ ),
    .B(\u_ppwm/u_ex/_312_ ),
    .A(\u_ppwm/u_ex/_310_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_735_  (.A1(\u_ppwm/u_ex/_310_ ),
    .A2(\u_ppwm/u_ex/_312_ ),
    .Y(\u_ppwm/u_ex/_314_ ),
    .B1(net315));
 sg13g2_a22oi_1 \u_ppwm/u_ex/_736_  (.Y(\u_ppwm/u_ex/_315_ ),
    .B1(net312),
    .B2(net385),
    .A2(net314),
    .A1(net383));
 sg13g2_nand3_1 \u_ppwm/u_ex/_737_  (.B(net307),
    .C(\u_ppwm/u_ex/_315_ ),
    .A(\u_ppwm/u_ex/_236_ ),
    .Y(\u_ppwm/u_ex/_316_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_738_  (.A1(\u_ppwm/u_ex/_313_ ),
    .A2(\u_ppwm/u_ex/_314_ ),
    .Y(\u_ppwm/u_ex/_317_ ),
    .B1(\u_ppwm/u_ex/_316_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_739_  (.B1(net439),
    .Y(\u_ppwm/u_ex/_318_ ),
    .A1(net384),
    .A2(net307));
 sg13g2_nor2_1 \u_ppwm/u_ex/_740_  (.A(\u_ppwm/u_ex/_317_ ),
    .B(\u_ppwm/u_ex/_318_ ),
    .Y(\u_ppwm/u_ex/_020_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_741_  (.Y(\u_ppwm/u_ex/_319_ ),
    .A(net383),
    .B(net322));
 sg13g2_nand3_1 \u_ppwm/u_ex/_742_  (.B(\u_ppwm/u_ex/_313_ ),
    .C(\u_ppwm/u_ex/_319_ ),
    .A(\u_ppwm/u_ex/_311_ ),
    .Y(\u_ppwm/u_ex/_320_ ));
 sg13g2_a21o_1 \u_ppwm/u_ex/_743_  (.A2(\u_ppwm/u_ex/_313_ ),
    .A1(\u_ppwm/u_ex/_311_ ),
    .B1(\u_ppwm/u_ex/_319_ ),
    .X(\u_ppwm/u_ex/_321_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_744_  (.B(\u_ppwm/u_ex/_320_ ),
    .C(\u_ppwm/u_ex/_321_ ),
    .A(net316),
    .Y(\u_ppwm/u_ex/_322_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_745_  (.B2(net658),
    .C1(\u_ppwm/u_ex/_295_ ),
    .B1(net312),
    .A1(net382),
    .Y(\u_ppwm/u_ex/_323_ ),
    .A2(net314));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_746_  (.B1(net441),
    .Y(\u_ppwm/u_ex/_324_ ),
    .A1(net383),
    .A2(net307));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_747_  (.A1(\u_ppwm/u_ex/_322_ ),
    .A2(\u_ppwm/u_ex/_323_ ),
    .Y(\u_ppwm/u_ex/_021_ ),
    .B1(\u_ppwm/u_ex/_324_ ));
 sg13g2_or2_1 \u_ppwm/u_ex/_748_  (.X(\u_ppwm/u_ex/_325_ ),
    .B(\u_ppwm/u_ex/_319_ ),
    .A(\u_ppwm/u_ex/_312_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_749_  (.B1(net322),
    .Y(\u_ppwm/u_ex/_326_ ),
    .A1(\u_ppwm/u_ex/reg_value_q[3] ),
    .A2(\u_ppwm/u_ex/reg_value_q[2] ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_750_  (.B1(\u_ppwm/u_ex/_326_ ),
    .Y(\u_ppwm/u_ex/_327_ ),
    .A1(\u_ppwm/u_ex/_310_ ),
    .A2(\u_ppwm/u_ex/_325_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_751_  (.Y(\u_ppwm/u_ex/_328_ ),
    .A(net382),
    .B(net321));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_752_  (.Y(\u_ppwm/u_ex/_329_ ),
    .A(net382),
    .B(net321));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_753_  (.Y(\u_ppwm/u_ex/_330_ ),
    .B(\u_ppwm/u_ex/_327_ ),
    .A_N(\u_ppwm/u_ex/_329_ ));
 sg13g2_nand2b_1 \u_ppwm/u_ex/_754_  (.Y(\u_ppwm/u_ex/_331_ ),
    .B(\u_ppwm/u_ex/_329_ ),
    .A_N(\u_ppwm/u_ex/_327_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_755_  (.B(\u_ppwm/u_ex/_330_ ),
    .C(\u_ppwm/u_ex/_331_ ),
    .A(net316),
    .Y(\u_ppwm/u_ex/_332_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_756_  (.B2(\u_ppwm/u_ex/reg_value_q[3] ),
    .C1(\u_ppwm/u_ex/_295_ ),
    .B1(net312),
    .A1(net381),
    .Y(\u_ppwm/u_ex/_333_ ),
    .A2(net314));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_757_  (.B1(net441),
    .Y(\u_ppwm/u_ex/_334_ ),
    .A1(net636),
    .A2(net307));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_758_  (.A1(\u_ppwm/u_ex/_332_ ),
    .A2(\u_ppwm/u_ex/_333_ ),
    .Y(\u_ppwm/u_ex/_022_ ),
    .B1(\u_ppwm/u_ex/_334_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_759_  (.Y(\u_ppwm/u_ex/_335_ ),
    .A(net381),
    .B(net321));
 sg13g2_a21o_1 \u_ppwm/u_ex/_760_  (.A2(\u_ppwm/u_ex/_330_ ),
    .A1(\u_ppwm/u_ex/_328_ ),
    .B1(\u_ppwm/u_ex/_335_ ),
    .X(\u_ppwm/u_ex/_336_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_761_  (.B(\u_ppwm/u_ex/_330_ ),
    .C(\u_ppwm/u_ex/_335_ ),
    .A(\u_ppwm/u_ex/_328_ ),
    .Y(\u_ppwm/u_ex/_337_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_762_  (.B(\u_ppwm/u_ex/_336_ ),
    .C(\u_ppwm/u_ex/_337_ ),
    .A(\u_ppwm/u_ex/_216_ ),
    .Y(\u_ppwm/u_ex/_338_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_763_  (.B2(net636),
    .C1(\u_ppwm/u_ex/_295_ ),
    .B1(\u_ppwm/u_ex/_227_ ),
    .A1(net380),
    .Y(\u_ppwm/u_ex/_339_ ),
    .A2(net314));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_764_  (.B1(net441),
    .Y(\u_ppwm/u_ex/_340_ ),
    .A1(net381),
    .A2(net307));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_765_  (.A1(\u_ppwm/u_ex/_338_ ),
    .A2(\u_ppwm/u_ex/_339_ ),
    .Y(\u_ppwm/u_ex/_023_ ),
    .B1(\u_ppwm/u_ex/_340_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_766_  (.Y(\u_ppwm/u_ex/_341_ ),
    .A(net380),
    .B(net321));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_767_  (.Y(\u_ppwm/u_ex/_342_ ),
    .A(net380),
    .B(net321));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_768_  (.B1(net321),
    .Y(\u_ppwm/u_ex/_343_ ),
    .A1(net381),
    .A2(\u_ppwm/u_ex/reg_value_q[4] ));
 sg13g2_inv_1 \u_ppwm/u_ex/_769_  (.Y(\u_ppwm/u_ex/_344_ ),
    .A(\u_ppwm/u_ex/_343_ ));
 sg13g2_nor2_1 \u_ppwm/u_ex/_770_  (.A(\u_ppwm/u_ex/_329_ ),
    .B(\u_ppwm/u_ex/_335_ ),
    .Y(\u_ppwm/u_ex/_345_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_771_  (.A1(\u_ppwm/u_ex/_327_ ),
    .A2(\u_ppwm/u_ex/_345_ ),
    .Y(\u_ppwm/u_ex/_346_ ),
    .B1(\u_ppwm/u_ex/_344_ ));
 sg13g2_or2_1 \u_ppwm/u_ex/_772_  (.X(\u_ppwm/u_ex/_347_ ),
    .B(\u_ppwm/u_ex/_346_ ),
    .A(\u_ppwm/u_ex/_342_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_773_  (.A1(\u_ppwm/u_ex/_342_ ),
    .A2(\u_ppwm/u_ex/_346_ ),
    .Y(\u_ppwm/u_ex/_348_ ),
    .B1(net315));
 sg13g2_nand2_1 \u_ppwm/u_ex/_774_  (.Y(\u_ppwm/u_ex/_349_ ),
    .A(\u_ppwm/u_ex/_347_ ),
    .B(\u_ppwm/u_ex/_348_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_775_  (.B2(\u_ppwm/u_ex/reg_value_q[5] ),
    .C1(\u_ppwm/u_ex/_295_ ),
    .B1(\u_ppwm/u_ex/_227_ ),
    .A1(\u_ppwm/u_ex/reg_value_q[7] ),
    .Y(\u_ppwm/u_ex/_350_ ),
    .A2(\u_ppwm/u_ex/_221_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_776_  (.B1(net441),
    .Y(\u_ppwm/u_ex/_351_ ),
    .A1(net639),
    .A2(net308));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_777_  (.A1(\u_ppwm/u_ex/_349_ ),
    .A2(\u_ppwm/u_ex/_350_ ),
    .Y(\u_ppwm/u_ex/_024_ ),
    .B1(\u_ppwm/u_ex/_351_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_778_  (.Y(\u_ppwm/u_ex/_352_ ),
    .A(\u_ppwm/u_ex/reg_value_q[7] ),
    .B(net321));
 sg13g2_nand3_1 \u_ppwm/u_ex/_779_  (.B(\u_ppwm/u_ex/_347_ ),
    .C(\u_ppwm/u_ex/_352_ ),
    .A(\u_ppwm/u_ex/_341_ ),
    .Y(\u_ppwm/u_ex/_353_ ));
 sg13g2_a21o_1 \u_ppwm/u_ex/_780_  (.A2(\u_ppwm/u_ex/_347_ ),
    .A1(\u_ppwm/u_ex/_341_ ),
    .B1(\u_ppwm/u_ex/_352_ ),
    .X(\u_ppwm/u_ex/_354_ ));
 sg13g2_nand3_1 \u_ppwm/u_ex/_781_  (.B(\u_ppwm/u_ex/_353_ ),
    .C(\u_ppwm/u_ex/_354_ ),
    .A(\u_ppwm/u_ex/_216_ ),
    .Y(\u_ppwm/u_ex/_355_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_782_  (.B2(net639),
    .C1(\u_ppwm/u_ex/_295_ ),
    .B1(\u_ppwm/u_ex/_227_ ),
    .A1(net379),
    .Y(\u_ppwm/u_ex/_356_ ),
    .A2(\u_ppwm/u_ex/_221_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_783_  (.B1(net441),
    .Y(\u_ppwm/u_ex/_357_ ),
    .A1(net653),
    .A2(net308));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_784_  (.A1(\u_ppwm/u_ex/_355_ ),
    .A2(\u_ppwm/u_ex/_356_ ),
    .Y(\u_ppwm/u_ex/_025_ ),
    .B1(\u_ppwm/u_ex/_357_ ));
 sg13g2_nor4_1 \u_ppwm/u_ex/_785_  (.A(\u_ppwm/u_ex/_329_ ),
    .B(\u_ppwm/u_ex/_335_ ),
    .C(\u_ppwm/u_ex/_342_ ),
    .D(\u_ppwm/u_ex/_352_ ),
    .Y(\u_ppwm/u_ex/_358_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_786_  (.B1(net321),
    .Y(\u_ppwm/u_ex/_359_ ),
    .A1(\u_ppwm/u_ex/reg_value_q[7] ),
    .A2(\u_ppwm/u_ex/reg_value_q[6] ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_787_  (.Y(\u_ppwm/u_ex/_360_ ),
    .A(\u_ppwm/u_ex/_343_ ),
    .B(\u_ppwm/u_ex/_359_ ));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_788_  (.A1(\u_ppwm/u_ex/_327_ ),
    .A2(\u_ppwm/u_ex/_358_ ),
    .Y(\u_ppwm/u_ex/_361_ ),
    .B1(\u_ppwm/u_ex/_360_ ));
 sg13g2_nand2_1 \u_ppwm/u_ex/_789_  (.Y(\u_ppwm/u_ex/_362_ ),
    .A(net379),
    .B(net322));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_790_  (.Y(\u_ppwm/u_ex/_363_ ),
    .A(net646),
    .B(net322));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_791_  (.A1(\u_ppwm/u_ex/_361_ ),
    .A2(\u_ppwm/u_ex/_363_ ),
    .Y(\u_ppwm/u_ex/_364_ ),
    .B1(\u_ppwm/u_ex/_217_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_792_  (.B1(\u_ppwm/u_ex/_364_ ),
    .Y(\u_ppwm/u_ex/_365_ ),
    .A1(\u_ppwm/u_ex/_361_ ),
    .A2(\u_ppwm/u_ex/_363_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_793_  (.B2(\u_ppwm/u_ex/reg_value_q[7] ),
    .C1(\u_ppwm/u_ex/_295_ ),
    .B1(net312),
    .A1(net378),
    .Y(\u_ppwm/u_ex/_366_ ),
    .A2(\u_ppwm/u_ex/_221_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_794_  (.B1(net441),
    .Y(\u_ppwm/u_ex/_367_ ),
    .A1(net646),
    .A2(net308));
 sg13g2_a21oi_1 \u_ppwm/u_ex/_795_  (.A1(\u_ppwm/u_ex/_365_ ),
    .A2(\u_ppwm/u_ex/_366_ ),
    .Y(\u_ppwm/u_ex/_026_ ),
    .B1(\u_ppwm/u_ex/_367_ ));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_796_  (.B1(\u_ppwm/u_ex/_362_ ),
    .Y(\u_ppwm/u_ex/_368_ ),
    .A1(\u_ppwm/u_ex/_361_ ),
    .A2(\u_ppwm/u_ex/_363_ ));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_797_  (.Y(\u_ppwm/u_ex/_369_ ),
    .A(net378),
    .B(net322));
 sg13g2_xnor2_1 \u_ppwm/u_ex/_798_  (.Y(\u_ppwm/u_ex/_370_ ),
    .A(\u_ppwm/u_ex/_368_ ),
    .B(\u_ppwm/u_ex/_369_ ));
 sg13g2_a221oi_1 \u_ppwm/u_ex/_799_  (.B2(\u_ppwm/u_ex/_216_ ),
    .C1(\u_ppwm/u_ex/_295_ ),
    .B1(\u_ppwm/u_ex/_370_ ),
    .A1(net646),
    .Y(\u_ppwm/u_ex/_371_ ),
    .A2(net312));
 sg13g2_o21ai_1 \u_ppwm/u_ex/_800_  (.B1(net441),
    .Y(\u_ppwm/u_ex/_372_ ),
    .A1(net378),
    .A2(net308));
 sg13g2_nor2_1 \u_ppwm/u_ex/_801_  (.A(\u_ppwm/u_ex/_371_ ),
    .B(\u_ppwm/u_ex/_372_ ),
    .Y(\u_ppwm/u_ex/_027_ ));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_802_  (.RESET_B(net51),
    .D(\u_ppwm/u_ex/_003_ ),
    .Q(\u_ppwm/pc[0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_803_  (.RESET_B(net44),
    .D(\u_ppwm/u_ex/_004_ ),
    .Q(\u_ppwm/pc[1] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_804_  (.RESET_B(net42),
    .D(\u_ppwm/u_ex/_005_ ),
    .Q(\u_ppwm/pc[2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_805_  (.RESET_B(net40),
    .D(net633),
    .Q(\u_ppwm/pc[3] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_806_  (.RESET_B(net38),
    .D(net629),
    .Q(\u_ppwm/u_ex/cmp_flag_q ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_807_  (.RESET_B(net36),
    .D(net650),
    .Q(\u_ppwm/pwm_value[0] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_808_  (.RESET_B(net34),
    .D(\u_ppwm/u_ex/_009_ ),
    .Q(\u_ppwm/pwm_value[1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_809_  (.RESET_B(net32),
    .D(\u_ppwm/u_ex/_010_ ),
    .Q(\u_ppwm/pwm_value[2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_810_  (.RESET_B(net30),
    .D(net665),
    .Q(\u_ppwm/pwm_value[3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_811_  (.RESET_B(net28),
    .D(net667),
    .Q(\u_ppwm/pwm_value[4] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_812_  (.RESET_B(net26),
    .D(\u_ppwm/u_ex/_013_ ),
    .Q(\u_ppwm/pwm_value[5] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_813_  (.RESET_B(net49),
    .D(net669),
    .Q(\u_ppwm/pwm_value[6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_814_  (.RESET_B(net47),
    .D(net674),
    .Q(\u_ppwm/pwm_value[7] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_815_  (.RESET_B(net45),
    .D(\u_ppwm/u_ex/_016_ ),
    .Q(\u_ppwm/pwm_value[8] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_816_  (.RESET_B(net41),
    .D(net652),
    .Q(\u_ppwm/pwm_value[9] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_817_  (.RESET_B(net37),
    .D(net635),
    .Q(\u_ppwm/u_ex/reg_value_q[0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_818_  (.RESET_B(net33),
    .D(net642),
    .Q(\u_ppwm/u_ex/reg_value_q[1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_819_  (.RESET_B(net29),
    .D(\u_ppwm/u_ex/_020_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_820_  (.RESET_B(net50),
    .D(net659),
    .Q(\u_ppwm/u_ex/reg_value_q[3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_821_  (.RESET_B(net46),
    .D(net637),
    .Q(\u_ppwm/u_ex/reg_value_q[4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_822_  (.RESET_B(net39),
    .D(\u_ppwm/u_ex/_023_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[5] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_823_  (.RESET_B(net31),
    .D(net640),
    .Q(\u_ppwm/u_ex/reg_value_q[6] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_824_  (.RESET_B(net48),
    .D(\u_ppwm/u_ex/_025_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[7] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_825_  (.RESET_B(net35),
    .D(net647),
    .Q(\u_ppwm/u_ex/reg_value_q[8] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_826_  (.RESET_B(net52),
    .D(\u_ppwm/u_ex/_027_ ),
    .Q(\u_ppwm/u_ex/reg_value_q[9] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_827_  (.RESET_B(net53),
    .D(net573),
    .Q(\u_ppwm/u_ex/state_q[0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_ex/_828_  (.RESET_B(net27),
    .D(\u_ppwm/u_ex/_001_ ),
    .Q(\u_ppwm/u_ex/state_q[1] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_ex/_829_  (.RESET_B(net43),
    .D(\u_ppwm/u_ex/_002_ ),
    .Q(\u_ppwm/u_ex/state_q[2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_tiehi \u_ppwm/u_ex/_828__27  (.L_HI(net27));
 sg13g2_tiehi \u_ppwm/u_ex/_811__28  (.L_HI(net28));
 sg13g2_tiehi \u_ppwm/u_ex/_819__29  (.L_HI(net29));
 sg13g2_tiehi \u_ppwm/u_ex/_810__30  (.L_HI(net30));
 sg13g2_tiehi \u_ppwm/u_ex/_823__31  (.L_HI(net31));
 sg13g2_tiehi \u_ppwm/u_ex/_809__32  (.L_HI(net32));
 sg13g2_tiehi \u_ppwm/u_ex/_818__33  (.L_HI(net33));
 sg13g2_tiehi \u_ppwm/u_ex/_808__34  (.L_HI(net34));
 sg13g2_tiehi \u_ppwm/u_ex/_825__35  (.L_HI(net35));
 sg13g2_tiehi \u_ppwm/u_ex/_807__36  (.L_HI(net36));
 sg13g2_tiehi \u_ppwm/u_ex/_817__37  (.L_HI(net37));
 sg13g2_tiehi \u_ppwm/u_ex/_806__38  (.L_HI(net38));
 sg13g2_tiehi \u_ppwm/u_ex/_822__39  (.L_HI(net39));
 sg13g2_tiehi \u_ppwm/u_ex/_805__40  (.L_HI(net40));
 sg13g2_tiehi \u_ppwm/u_ex/_816__41  (.L_HI(net41));
 sg13g2_tiehi \u_ppwm/u_ex/_804__42  (.L_HI(net42));
 sg13g2_tiehi \u_ppwm/u_ex/_829__43  (.L_HI(net43));
 sg13g2_tiehi \u_ppwm/u_ex/_803__44  (.L_HI(net44));
 sg13g2_tiehi \u_ppwm/u_ex/_815__45  (.L_HI(net45));
 sg13g2_tiehi \u_ppwm/u_ex/_821__46  (.L_HI(net46));
 sg13g2_tiehi \u_ppwm/u_ex/_814__47  (.L_HI(net47));
 sg13g2_tiehi \u_ppwm/u_ex/_824__48  (.L_HI(net48));
 sg13g2_tiehi \u_ppwm/u_ex/_813__49  (.L_HI(net49));
 sg13g2_tiehi \u_ppwm/u_ex/_820__50  (.L_HI(net50));
 sg13g2_tiehi \u_ppwm/u_ex/_802__51  (.L_HI(net51));
 sg13g2_tiehi \u_ppwm/u_ex/_826__52  (.L_HI(net52));
 sg13g2_tiehi \u_ppwm/u_ex/_827__53  (.L_HI(net53));
 sg13g2_tiehi \u_ppwm/u_mem/_1190__54  (.L_HI(net54));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_053_  (.Y(\u_ppwm/u_global_counter/_020_ ),
    .A(net546));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_054_  (.Y(\u_ppwm/u_global_counter/_021_ ),
    .A(net609));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_055_  (.Y(\u_ppwm/u_global_counter/_022_ ),
    .A(net615));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_056_  (.Y(\u_ppwm/u_global_counter/_023_ ),
    .A(net577));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_057_  (.Y(\u_ppwm/u_global_counter/_024_ ),
    .A(net614));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_058_  (.Y(\u_ppwm/u_global_counter/_025_ ),
    .A(net564));
 sg13g2_inv_1 \u_ppwm/u_global_counter/_059_  (.Y(\u_ppwm/u_global_counter/_026_ ),
    .A(net336));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_060_  (.B(net336),
    .A(net268),
    .X(\u_ppwm/u_global_counter/_000_ ));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_061_  (.B(net654),
    .C(net336),
    .A(net268),
    .Y(\u_ppwm/u_global_counter/_027_ ));
 sg13g2_a21o_1 \u_ppwm/u_global_counter/_062_  (.A2(net336),
    .A1(net268),
    .B1(net654),
    .X(\u_ppwm/u_global_counter/_028_ ));
 sg13g2_and2_1 \u_ppwm/u_global_counter/_063_  (.A(\u_ppwm/u_global_counter/_027_ ),
    .B(net655),
    .X(\u_ppwm/u_global_counter/_001_ ));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_064_  (.B(\u_ppwm/global_counter_high[1] ),
    .C(net251),
    .A(net268),
    .Y(\u_ppwm/u_global_counter/_029_ ),
    .D(net336));
 sg13g2_xnor2_1 \u_ppwm/u_global_counter/_065_  (.Y(\u_ppwm/u_global_counter/_002_ ),
    .A(net251),
    .B(\u_ppwm/u_global_counter/_027_ ));
 sg13g2_nor2_1 \u_ppwm/u_global_counter/_066_  (.A(\u_ppwm/u_global_counter/_020_ ),
    .B(\u_ppwm/u_global_counter/_029_ ),
    .Y(\u_ppwm/u_global_counter/_030_ ));
 sg13g2_xnor2_1 \u_ppwm/u_global_counter/_067_  (.Y(\u_ppwm/u_global_counter/_003_ ),
    .A(net546),
    .B(\u_ppwm/u_global_counter/_029_ ));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_068_  (.B(\u_ppwm/u_global_counter/_030_ ),
    .A(net528),
    .X(\u_ppwm/u_global_counter/_004_ ));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_069_  (.B(net546),
    .C(net528),
    .A(net251),
    .Y(\u_ppwm/u_global_counter/_031_ ),
    .D(net586));
 sg13g2_nor2_1 \u_ppwm/u_global_counter/_070_  (.A(\u_ppwm/u_global_counter/_027_ ),
    .B(\u_ppwm/u_global_counter/_031_ ),
    .Y(\u_ppwm/u_global_counter/_032_ ));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_071_  (.A1(net528),
    .A2(\u_ppwm/u_global_counter/_030_ ),
    .Y(\u_ppwm/u_global_counter/_033_ ),
    .B1(net586));
 sg13g2_nor2_1 \u_ppwm/u_global_counter/_072_  (.A(\u_ppwm/u_global_counter/_032_ ),
    .B(net587),
    .Y(\u_ppwm/u_global_counter/_005_ ));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_073_  (.B(\u_ppwm/u_global_counter/_032_ ),
    .A(net202),
    .X(\u_ppwm/u_global_counter/_006_ ));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_074_  (.B(\u_ppwm/global_counter_high[1] ),
    .C(net202),
    .A(net268),
    .Y(\u_ppwm/u_global_counter/_034_ ),
    .D(net461));
 sg13g2_nor3_2 \u_ppwm/u_global_counter/_075_  (.A(\u_ppwm/u_global_counter/_026_ ),
    .B(\u_ppwm/u_global_counter/_031_ ),
    .C(\u_ppwm/u_global_counter/_034_ ),
    .Y(\u_ppwm/u_global_counter/_035_ ));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_076_  (.A1(net202),
    .A2(\u_ppwm/u_global_counter/_032_ ),
    .Y(\u_ppwm/u_global_counter/_036_ ),
    .B1(net461));
 sg13g2_nor2_1 \u_ppwm/u_global_counter/_077_  (.A(\u_ppwm/u_global_counter/_035_ ),
    .B(net462),
    .Y(\u_ppwm/u_global_counter/_007_ ));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_078_  (.B(\u_ppwm/u_global_counter/_035_ ),
    .A(net291),
    .X(\u_ppwm/u_global_counter/_008_ ));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_079_  (.B(net657),
    .C(\u_ppwm/u_global_counter/_035_ ),
    .A(net291),
    .Y(\u_ppwm/u_global_counter/_037_ ));
 sg13g2_a21o_1 \u_ppwm/u_global_counter/_080_  (.A2(\u_ppwm/u_global_counter/_035_ ),
    .A1(net291),
    .B1(net657),
    .X(\u_ppwm/u_global_counter/_038_ ));
 sg13g2_and2_1 \u_ppwm/u_global_counter/_081_  (.A(\u_ppwm/u_global_counter/_037_ ),
    .B(\u_ppwm/u_global_counter/_038_ ),
    .X(\u_ppwm/u_global_counter/_009_ ));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_082_  (.B(\u_ppwm/global_counter_high[9] ),
    .C(net227),
    .A(net291),
    .Y(\u_ppwm/u_global_counter/_039_ ),
    .D(\u_ppwm/u_global_counter/_035_ ));
 sg13g2_xnor2_1 \u_ppwm/u_global_counter/_083_  (.Y(\u_ppwm/u_global_counter/_010_ ),
    .A(net227),
    .B(\u_ppwm/u_global_counter/_037_ ));
 sg13g2_nand4_1 \u_ppwm/u_global_counter/_084_  (.B(\u_ppwm/global_counter_high[9] ),
    .C(net227),
    .A(net291),
    .Y(\u_ppwm/u_global_counter/_040_ ),
    .D(net609));
 sg13g2_nor3_2 \u_ppwm/u_global_counter/_085_  (.A(\u_ppwm/u_global_counter/_031_ ),
    .B(\u_ppwm/u_global_counter/_034_ ),
    .C(\u_ppwm/u_global_counter/_040_ ),
    .Y(\u_ppwm/u_global_counter/_041_ ));
 sg13g2_a22oi_1 \u_ppwm/u_global_counter/_086_  (.Y(\u_ppwm/u_global_counter/_011_ ),
    .B1(\u_ppwm/u_global_counter/_041_ ),
    .B2(net336),
    .A2(\u_ppwm/u_global_counter/_039_ ),
    .A1(\u_ppwm/u_global_counter/_021_ ));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_087_  (.A1(\u_ppwm/period_start ),
    .A2(net331),
    .Y(\u_ppwm/u_global_counter/_042_ ),
    .B1(net555));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_088_  (.B(\u_ppwm/period_start ),
    .C(net331),
    .A(net555),
    .Y(\u_ppwm/u_global_counter/_043_ ));
 sg13g2_nor2b_1 \u_ppwm/u_global_counter/_089_  (.A(net556),
    .B_N(\u_ppwm/u_global_counter/_043_ ),
    .Y(\u_ppwm/u_global_counter/_012_ ));
 sg13g2_and3_2 \u_ppwm/u_global_counter/_090_  (.X(\u_ppwm/u_global_counter/_044_ ),
    .A(net555),
    .B(net615),
    .C(\u_ppwm/period_start ));
 sg13g2_a22oi_1 \u_ppwm/u_global_counter/_091_  (.Y(\u_ppwm/u_global_counter/_013_ ),
    .B1(\u_ppwm/u_global_counter/_044_ ),
    .B2(net331),
    .A2(\u_ppwm/u_global_counter/_043_ ),
    .A1(\u_ppwm/u_global_counter/_022_ ));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_092_  (.A1(net331),
    .A2(\u_ppwm/u_global_counter/_044_ ),
    .Y(\u_ppwm/u_global_counter/_045_ ),
    .B1(net552));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_093_  (.B(net331),
    .C(\u_ppwm/u_global_counter/_044_ ),
    .A(net552),
    .Y(\u_ppwm/u_global_counter/_046_ ));
 sg13g2_nor2b_1 \u_ppwm/u_global_counter/_094_  (.A(net553),
    .B_N(\u_ppwm/u_global_counter/_046_ ),
    .Y(\u_ppwm/u_global_counter/_014_ ));
 sg13g2_and3_2 \u_ppwm/u_global_counter/_095_  (.X(\u_ppwm/u_global_counter/_047_ ),
    .A(net552),
    .B(net577),
    .C(\u_ppwm/u_global_counter/_044_ ));
 sg13g2_and2_1 \u_ppwm/u_global_counter/_096_  (.A(net331),
    .B(\u_ppwm/u_global_counter/_047_ ),
    .X(\u_ppwm/u_global_counter/_048_ ));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_097_  (.A1(\u_ppwm/u_global_counter/_023_ ),
    .A2(\u_ppwm/u_global_counter/_046_ ),
    .Y(\u_ppwm/u_global_counter/_015_ ),
    .B1(\u_ppwm/u_global_counter/_048_ ));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_098_  (.B(net331),
    .C(\u_ppwm/u_global_counter/_047_ ),
    .A(net198),
    .Y(\u_ppwm/u_global_counter/_049_ ));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_099_  (.B(\u_ppwm/u_global_counter/_048_ ),
    .A(net198),
    .X(\u_ppwm/u_global_counter/_016_ ));
 sg13g2_and2_1 \u_ppwm/u_global_counter/_100_  (.A(net198),
    .B(net614),
    .X(\u_ppwm/u_global_counter/_050_ ));
 sg13g2_nand3_1 \u_ppwm/u_global_counter/_101_  (.B(\u_ppwm/u_global_counter/_047_ ),
    .C(\u_ppwm/u_global_counter/_050_ ),
    .A(\u_ppwm/u_global_counter/_041_ ),
    .Y(\u_ppwm/u_global_counter/_051_ ));
 sg13g2_a22oi_1 \u_ppwm/u_global_counter/_102_  (.Y(\u_ppwm/u_global_counter/_017_ ),
    .B1(\u_ppwm/u_global_counter/_050_ ),
    .B2(\u_ppwm/u_global_counter/_048_ ),
    .A2(\u_ppwm/u_global_counter/_049_ ),
    .A1(\u_ppwm/u_global_counter/_024_ ));
 sg13g2_and4_1 \u_ppwm/u_global_counter/_103_  (.A(net564),
    .B(net331),
    .C(\u_ppwm/u_global_counter/_047_ ),
    .D(\u_ppwm/u_global_counter/_050_ ),
    .X(\u_ppwm/u_global_counter/_052_ ));
 sg13g2_a21oi_1 \u_ppwm/u_global_counter/_104_  (.A1(\u_ppwm/u_global_counter/_025_ ),
    .A2(\u_ppwm/u_global_counter/_051_ ),
    .Y(\u_ppwm/u_global_counter/_018_ ),
    .B1(\u_ppwm/u_global_counter/_052_ ));
 sg13g2_xor2_1 \u_ppwm/u_global_counter/_105_  (.B(\u_ppwm/u_global_counter/_052_ ),
    .A(net204),
    .X(\u_ppwm/u_global_counter/_019_ ));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_106_  (.RESET_B(net438),
    .D(net269),
    .Q(\u_ppwm/global_counter_high[0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_107_  (.RESET_B(net438),
    .D(net656),
    .Q(\u_ppwm/global_counter_high[1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_108_  (.RESET_B(net438),
    .D(net252),
    .Q(\u_ppwm/global_counter_high[2] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_109_  (.RESET_B(net438),
    .D(net547),
    .Q(\u_ppwm/global_counter_high[3] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_110_  (.RESET_B(net440),
    .D(net529),
    .Q(\u_ppwm/global_counter_high[4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_111_  (.RESET_B(net438),
    .D(net588),
    .Q(\u_ppwm/global_counter_high[5] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_112_  (.RESET_B(net439),
    .D(net203),
    .Q(\u_ppwm/global_counter_high[6] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_113_  (.RESET_B(net438),
    .D(net463),
    .Q(\u_ppwm/global_counter_high[7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_114_  (.RESET_B(net439),
    .D(net292),
    .Q(\u_ppwm/global_counter_high[8] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_115_  (.RESET_B(net439),
    .D(\u_ppwm/u_global_counter/_009_ ),
    .Q(\u_ppwm/global_counter_high[9] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_116_  (.RESET_B(net438),
    .D(net228),
    .Q(\u_ppwm/global_counter_high[10] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_117_  (.RESET_B(net438),
    .D(net610),
    .Q(\u_ppwm/global_counter_high[11] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_118_  (.RESET_B(net440),
    .D(net557),
    .Q(\u_ppwm/global_counter_high[12] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_119_  (.RESET_B(net440),
    .D(net616),
    .Q(\u_ppwm/global_counter_high[13] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_120_  (.RESET_B(net440),
    .D(net554),
    .Q(\u_ppwm/global_counter_high[14] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_121_  (.RESET_B(net440),
    .D(net578),
    .Q(\u_ppwm/global_counter_high[15] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_122_  (.RESET_B(net440),
    .D(net199),
    .Q(\u_ppwm/global_counter_high[16] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_123_  (.RESET_B(net440),
    .D(\u_ppwm/u_global_counter/_017_ ),
    .Q(\u_ppwm/global_counter_high[17] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_124_  (.RESET_B(net440),
    .D(net565),
    .Q(\u_ppwm/global_counter_high[18] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_global_counter/_125_  (.RESET_B(net441),
    .D(net205),
    .Q(\u_ppwm/global_counter_high[19] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_inv_1 \u_ppwm/u_mem/_0613_  (.Y(\u_ppwm/u_mem/_0126_ ),
    .A(net206));
 sg13g2_inv_1 \u_ppwm/u_mem/_0614_  (.Y(\u_ppwm/u_mem/_0127_ ),
    .A(net1));
 sg13g2_inv_1 \u_ppwm/u_mem/_0615_  (.Y(\u_ppwm/u_mem/_0128_ ),
    .A(net521));
 sg13g2_inv_1 \u_ppwm/u_mem/_0616_  (.Y(\u_ppwm/u_mem/_0129_ ),
    .A(net592));
 sg13g2_inv_1 \u_ppwm/u_mem/_0617_  (.Y(\u_ppwm/u_mem/_0130_ ),
    .A(net558));
 sg13g2_inv_1 \u_ppwm/u_mem/_0618_  (.Y(\u_ppwm/u_mem/_0131_ ),
    .A(net543));
 sg13g2_inv_1 \u_ppwm/u_mem/_0619_  (.Y(\u_ppwm/u_mem/_0132_ ),
    .A(net233));
 sg13g2_inv_1 \u_ppwm/u_mem/_0620_  (.Y(\u_ppwm/u_mem/_0133_ ),
    .A(net566));
 sg13g2_inv_1 \u_ppwm/u_mem/_0621_  (.Y(\u_ppwm/u_mem/_0134_ ),
    .A(net477));
 sg13g2_inv_1 \u_ppwm/u_mem/_0622_  (.Y(\u_ppwm/u_mem/_0135_ ),
    .A(net534));
 sg13g2_inv_1 \u_ppwm/u_mem/_0623_  (.Y(\u_ppwm/u_mem/_0136_ ),
    .A(net471));
 sg13g2_inv_1 \u_ppwm/u_mem/_0624_  (.Y(\u_ppwm/u_mem/_0137_ ),
    .A(net579));
 sg13g2_inv_1 \u_ppwm/u_mem/_0625_  (.Y(\u_ppwm/u_mem/_0138_ ),
    .A(net286));
 sg13g2_inv_1 \u_ppwm/u_mem/_0626_  (.Y(\u_ppwm/u_mem/_0139_ ),
    .A(net212));
 sg13g2_inv_1 \u_ppwm/u_mem/_0627_  (.Y(\u_ppwm/u_mem/_0140_ ),
    .A(net262));
 sg13g2_inv_1 \u_ppwm/u_mem/_0628_  (.Y(\u_ppwm/u_mem/_0141_ ),
    .A(net489));
 sg13g2_inv_1 \u_ppwm/u_mem/_0629_  (.Y(\u_ppwm/u_mem/_0142_ ),
    .A(net473));
 sg13g2_inv_1 \u_ppwm/u_mem/_0630_  (.Y(\u_ppwm/u_mem/_0143_ ),
    .A(net295));
 sg13g2_inv_1 \u_ppwm/u_mem/_0631_  (.Y(\u_ppwm/u_mem/_0144_ ),
    .A(net458));
 sg13g2_inv_1 \u_ppwm/u_mem/_0632_  (.Y(\u_ppwm/u_mem/_0145_ ),
    .A(net274));
 sg13g2_inv_1 \u_ppwm/u_mem/_0633_  (.Y(\u_ppwm/u_mem/_0146_ ),
    .A(net498));
 sg13g2_inv_1 \u_ppwm/u_mem/_0634_  (.Y(\u_ppwm/u_mem/_0147_ ),
    .A(net266));
 sg13g2_inv_1 \u_ppwm/u_mem/_0635_  (.Y(\u_ppwm/u_mem/_0148_ ),
    .A(net210));
 sg13g2_inv_1 \u_ppwm/u_mem/_0636_  (.Y(\u_ppwm/u_mem/_0149_ ),
    .A(net245));
 sg13g2_inv_1 \u_ppwm/u_mem/_0637_  (.Y(\u_ppwm/u_mem/_0150_ ),
    .A(net258));
 sg13g2_inv_1 \u_ppwm/u_mem/_0638_  (.Y(\u_ppwm/u_mem/_0151_ ),
    .A(net284));
 sg13g2_inv_1 \u_ppwm/u_mem/_0639_  (.Y(\u_ppwm/u_mem/_0152_ ),
    .A(net231));
 sg13g2_inv_1 \u_ppwm/u_mem/_0640_  (.Y(\u_ppwm/u_mem/_0153_ ),
    .A(net485));
 sg13g2_inv_1 \u_ppwm/u_mem/_0641_  (.Y(\u_ppwm/u_mem/_0154_ ),
    .A(net574));
 sg13g2_inv_1 \u_ppwm/u_mem/_0642_  (.Y(\u_ppwm/u_mem/_0155_ ),
    .A(net516));
 sg13g2_inv_1 \u_ppwm/u_mem/_0643_  (.Y(\u_ppwm/u_mem/_0156_ ),
    .A(net225));
 sg13g2_inv_1 \u_ppwm/u_mem/_0644_  (.Y(\u_ppwm/u_mem/_0157_ ),
    .A(net239));
 sg13g2_inv_1 \u_ppwm/u_mem/_0645_  (.Y(\u_ppwm/u_mem/_0158_ ),
    .A(net508));
 sg13g2_inv_1 \u_ppwm/u_mem/_0646_  (.Y(\u_ppwm/u_mem/_0159_ ),
    .A(net538));
 sg13g2_inv_1 \u_ppwm/u_mem/_0647_  (.Y(\u_ppwm/u_mem/_0160_ ),
    .A(net229));
 sg13g2_inv_1 \u_ppwm/u_mem/_0648_  (.Y(\u_ppwm/u_mem/_0161_ ),
    .A(net525));
 sg13g2_inv_1 \u_ppwm/u_mem/_0649_  (.Y(\u_ppwm/u_mem/_0162_ ),
    .A(net544));
 sg13g2_inv_1 \u_ppwm/u_mem/_0650_  (.Y(\u_ppwm/u_mem/_0163_ ),
    .A(net524));
 sg13g2_inv_1 \u_ppwm/u_mem/_0651_  (.Y(\u_ppwm/u_mem/_0164_ ),
    .A(net293));
 sg13g2_inv_1 \u_ppwm/u_mem/_0652_  (.Y(\u_ppwm/u_mem/_0165_ ),
    .A(net510));
 sg13g2_inv_1 \u_ppwm/u_mem/_0653_  (.Y(\u_ppwm/u_mem/_0166_ ),
    .A(net278));
 sg13g2_inv_1 \u_ppwm/u_mem/_0654_  (.Y(\u_ppwm/u_mem/_0167_ ),
    .A(net276));
 sg13g2_inv_1 \u_ppwm/u_mem/_0655_  (.Y(\u_ppwm/u_mem/_0168_ ),
    .A(net453));
 sg13g2_inv_1 \u_ppwm/u_mem/_0656_  (.Y(\u_ppwm/u_mem/_0169_ ),
    .A(net620));
 sg13g2_inv_1 \u_ppwm/u_mem/_0657_  (.Y(\u_ppwm/u_mem/_0170_ ),
    .A(net208));
 sg13g2_inv_1 \u_ppwm/u_mem/_0658_  (.Y(\u_ppwm/u_mem/_0171_ ),
    .A(net243));
 sg13g2_inv_1 \u_ppwm/u_mem/_0659_  (.Y(\u_ppwm/u_mem/_0172_ ),
    .A(net303));
 sg13g2_inv_1 \u_ppwm/u_mem/_0660_  (.Y(\u_ppwm/u_mem/_0173_ ),
    .A(net270));
 sg13g2_inv_1 \u_ppwm/u_mem/_0661_  (.Y(\u_ppwm/u_mem/_0174_ ),
    .A(net467));
 sg13g2_inv_1 \u_ppwm/u_mem/_0662_  (.Y(\u_ppwm/u_mem/_0175_ ),
    .A(net487));
 sg13g2_inv_1 \u_ppwm/u_mem/_0663_  (.Y(\u_ppwm/u_mem/_0176_ ),
    .A(net617));
 sg13g2_inv_1 \u_ppwm/u_mem/_0664_  (.Y(\u_ppwm/u_mem/_0177_ ),
    .A(net287));
 sg13g2_inv_1 \u_ppwm/u_mem/_0665_  (.Y(\u_ppwm/u_mem/_0178_ ),
    .A(net493));
 sg13g2_inv_1 \u_ppwm/u_mem/_0666_  (.Y(\u_ppwm/u_mem/_0179_ ),
    .A(net253));
 sg13g2_inv_1 \u_ppwm/u_mem/_0667_  (.Y(\u_ppwm/u_mem/_0180_ ),
    .A(net224));
 sg13g2_inv_1 \u_ppwm/u_mem/_0668_  (.Y(\u_ppwm/u_mem/_0181_ ),
    .A(net214));
 sg13g2_inv_1 \u_ppwm/u_mem/_0669_  (.Y(\u_ppwm/u_mem/_0182_ ),
    .A(net282));
 sg13g2_inv_1 \u_ppwm/u_mem/_0670_  (.Y(\u_ppwm/u_mem/_0183_ ),
    .A(net559));
 sg13g2_inv_1 \u_ppwm/u_mem/_0671_  (.Y(\u_ppwm/u_mem/_0184_ ),
    .A(net256));
 sg13g2_inv_1 \u_ppwm/u_mem/_0672_  (.Y(\u_ppwm/u_mem/_0185_ ),
    .A(net576));
 sg13g2_inv_1 \u_ppwm/u_mem/_0673_  (.Y(\u_ppwm/u_mem/_0186_ ),
    .A(net306));
 sg13g2_inv_1 \u_ppwm/u_mem/_0674_  (.Y(\u_ppwm/u_mem/_0187_ ),
    .A(net237));
 sg13g2_inv_1 \u_ppwm/u_mem/_0675_  (.Y(\u_ppwm/u_mem/_0188_ ),
    .A(net260));
 sg13g2_inv_1 \u_ppwm/u_mem/_0676_  (.Y(\u_ppwm/u_mem/_0189_ ),
    .A(net515));
 sg13g2_inv_1 \u_ppwm/u_mem/_0677_  (.Y(\u_ppwm/u_mem/_0190_ ),
    .A(net247));
 sg13g2_inv_1 \u_ppwm/u_mem/_0678_  (.Y(\u_ppwm/u_mem/_0191_ ),
    .A(net455));
 sg13g2_inv_1 \u_ppwm/u_mem/_0679_  (.Y(\u_ppwm/u_mem/_0192_ ),
    .A(net457));
 sg13g2_inv_1 \u_ppwm/u_mem/_0680_  (.Y(\u_ppwm/u_mem/_0193_ ),
    .A(net297));
 sg13g2_inv_1 \u_ppwm/u_mem/_0681_  (.Y(\u_ppwm/u_mem/_0194_ ),
    .A(net548));
 sg13g2_inv_1 \u_ppwm/u_mem/_0682_  (.Y(\u_ppwm/u_mem/_0195_ ),
    .A(net519));
 sg13g2_inv_1 \u_ppwm/u_mem/_0683_  (.Y(\u_ppwm/u_mem/_0196_ ),
    .A(net539));
 sg13g2_inv_1 \u_ppwm/u_mem/_0684_  (.Y(\u_ppwm/u_mem/_0197_ ),
    .A(net541));
 sg13g2_inv_1 \u_ppwm/u_mem/_0685_  (.Y(\u_ppwm/u_mem/_0198_ ),
    .A(net545));
 sg13g2_inv_1 \u_ppwm/u_mem/_0686_  (.Y(\u_ppwm/u_mem/_0199_ ),
    .A(net280));
 sg13g2_inv_1 \u_ppwm/u_mem/_0687_  (.Y(\u_ppwm/u_mem/_0200_ ),
    .A(net466));
 sg13g2_inv_1 \u_ppwm/u_mem/_0688_  (.Y(\u_ppwm/u_mem/_0201_ ),
    .A(net459));
 sg13g2_inv_1 \u_ppwm/u_mem/_0689_  (.Y(\u_ppwm/u_mem/_0202_ ),
    .A(net494));
 sg13g2_inv_1 \u_ppwm/u_mem/_0690_  (.Y(\u_ppwm/u_mem/_0203_ ),
    .A(net289));
 sg13g2_inv_1 \u_ppwm/u_mem/_0691_  (.Y(\u_ppwm/u_mem/_0204_ ),
    .A(net606));
 sg13g2_inv_1 \u_ppwm/u_mem/_0692_  (.Y(\u_ppwm/u_mem/_0205_ ),
    .A(net272));
 sg13g2_inv_1 \u_ppwm/u_mem/_0693_  (.Y(\u_ppwm/u_mem/_0206_ ),
    .A(net216));
 sg13g2_inv_1 \u_ppwm/u_mem/_0694_  (.Y(\u_ppwm/u_mem/_0207_ ),
    .A(net517));
 sg13g2_inv_1 \u_ppwm/u_mem/_0695_  (.Y(\u_ppwm/u_mem/_0208_ ),
    .A(net530));
 sg13g2_inv_1 \u_ppwm/u_mem/_0696_  (.Y(\u_ppwm/u_mem/_0209_ ),
    .A(net575));
 sg13g2_inv_1 \u_ppwm/u_mem/_0697_  (.Y(\u_ppwm/u_mem/_0210_ ),
    .A(net235));
 sg13g2_inv_1 \u_ppwm/u_mem/_0698_  (.Y(\u_ppwm/u_mem/_0211_ ),
    .A(net254));
 sg13g2_inv_1 \u_ppwm/u_mem/_0699_  (.Y(\u_ppwm/u_mem/_0212_ ),
    .A(net570));
 sg13g2_inv_1 \u_ppwm/u_mem/_0700_  (.Y(\u_ppwm/u_mem/_0213_ ),
    .A(net299));
 sg13g2_inv_1 \u_ppwm/u_mem/_0701_  (.Y(\u_ppwm/u_mem/_0214_ ),
    .A(net475));
 sg13g2_inv_1 \u_ppwm/u_mem/_0702_  (.Y(\u_ppwm/u_mem/_0215_ ),
    .A(net505));
 sg13g2_inv_1 \u_ppwm/u_mem/_0703_  (.Y(\u_ppwm/u_mem/_0216_ ),
    .A(net500));
 sg13g2_inv_1 \u_ppwm/u_mem/_0704_  (.Y(\u_ppwm/u_mem/_0217_ ),
    .A(net479));
 sg13g2_inv_1 \u_ppwm/u_mem/_0705_  (.Y(\u_ppwm/u_mem/_0218_ ),
    .A(net537));
 sg13g2_inv_1 \u_ppwm/u_mem/_0706_  (.Y(\u_ppwm/u_mem/_0219_ ),
    .A(net503));
 sg13g2_inv_1 \u_ppwm/u_mem/_0707_  (.Y(\u_ppwm/u_mem/_0220_ ),
    .A(net301));
 sg13g2_inv_1 \u_ppwm/u_mem/_0708_  (.Y(\u_ppwm/u_mem/_0221_ ),
    .A(net483));
 sg13g2_inv_1 \u_ppwm/u_mem/_0709_  (.Y(\u_ppwm/u_mem/_0222_ ),
    .A(net591));
 sg13g2_inv_1 \u_ppwm/u_mem/_0710_  (.Y(\u_ppwm/u_mem/_0223_ ),
    .A(net589));
 sg13g2_inv_1 \u_ppwm/u_mem/_0711_  (.Y(\u_ppwm/u_mem/_0224_ ),
    .A(net506));
 sg13g2_inv_1 \u_ppwm/u_mem/_0712_  (.Y(\u_ppwm/u_mem/_0225_ ),
    .A(net491));
 sg13g2_inv_1 \u_ppwm/u_mem/_0713_  (.Y(\u_ppwm/u_mem/_0226_ ),
    .A(net469));
 sg13g2_inv_1 \u_ppwm/u_mem/_0714_  (.Y(\u_ppwm/u_mem/_0227_ ),
    .A(net464));
 sg13g2_inv_1 \u_ppwm/u_mem/_0715_  (.Y(\u_ppwm/u_mem/_0228_ ),
    .A(net523));
 sg13g2_inv_1 \u_ppwm/u_mem/_0716_  (.Y(\u_ppwm/u_mem/_0229_ ),
    .A(net241));
 sg13g2_inv_1 \u_ppwm/u_mem/_0717_  (.Y(\u_ppwm/u_mem/_0230_ ),
    .A(net560));
 sg13g2_inv_1 \u_ppwm/u_mem/_0718_  (.Y(\u_ppwm/u_mem/_0231_ ),
    .A(net481));
 sg13g2_inv_1 \u_ppwm/u_mem/_0719_  (.Y(\u_ppwm/u_mem/_0232_ ),
    .A(net600));
 sg13g2_inv_1 \u_ppwm/u_mem/_0720_  (.Y(\u_ppwm/u_mem/_0233_ ),
    .A(net532));
 sg13g2_inv_1 \u_ppwm/u_mem/_0721_  (.Y(\u_ppwm/u_mem/_0234_ ),
    .A(net527));
 sg13g2_inv_1 \u_ppwm/u_mem/_0722_  (.Y(\u_ppwm/u_mem/_0235_ ),
    .A(net501));
 sg13g2_inv_1 \u_ppwm/u_mem/_0723_  (.Y(\u_ppwm/u_mem/_0236_ ),
    .A(net585));
 sg13g2_inv_1 \u_ppwm/u_mem/_0724_  (.Y(\u_ppwm/u_mem/_0237_ ),
    .A(net511));
 sg13g2_inv_2 \u_ppwm/u_mem/_0725_  (.Y(\u_ppwm/u_mem/_0238_ ),
    .A(net423));
 sg13g2_inv_1 \u_ppwm/u_mem/_0726_  (.Y(\u_ppwm/u_mem/_0239_ ),
    .A(net513));
 sg13g2_inv_1 \u_ppwm/u_mem/_0727_  (.Y(\u_ppwm/u_mem/_0240_ ),
    .A(net408));
 sg13g2_inv_2 \u_ppwm/u_mem/_0728_  (.Y(\u_ppwm/u_mem/_0241_ ),
    .A(net402));
 sg13g2_inv_4 \u_ppwm/u_mem/_0729_  (.A(net400),
    .Y(\u_ppwm/u_mem/_0242_ ));
 sg13g2_nor3_1 \u_ppwm/u_mem/_0730_  (.A(\u_ppwm/u_mem/_0127_ ),
    .B(\u_ppwm/u_mem/_0238_ ),
    .C(\u_ppwm/mem_write_done ),
    .Y(\u_ppwm/u_mem/_0243_ ));
 sg13g2_nor2_1 \u_ppwm/u_mem/_0731_  (.A(net1),
    .B(\u_ppwm/u_mem/_0238_ ),
    .Y(\u_ppwm/u_mem/_0244_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0732_  (.A1(\u_ppwm/u_mem/_0239_ ),
    .A2(\u_ppwm/u_mem/_0244_ ),
    .Y(\u_ppwm/u_mem/_0004_ ),
    .B1(\u_ppwm/u_mem/_0243_ ));
 sg13g2_nand3_1 \u_ppwm/u_mem/_0733_  (.B(net597),
    .C(net624),
    .A(net549),
    .Y(\u_ppwm/u_mem/_0245_ ));
 sg13g2_nand3_1 \u_ppwm/u_mem/_0734_  (.B(net619),
    .C(net618),
    .A(net582),
    .Y(\u_ppwm/u_mem/_0246_ ));
 sg13g2_nor3_1 \u_ppwm/u_mem/_0735_  (.A(net602),
    .B(\u_ppwm/u_mem/_0245_ ),
    .C(\u_ppwm/u_mem/_0246_ ),
    .Y(\u_ppwm/u_mem/_0247_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0736_  (.Y(\u_ppwm/u_mem/_0248_ ),
    .A(net338),
    .B(net423));
 sg13g2_nor4_1 \u_ppwm/u_mem/_0737_  (.A(net602),
    .B(\u_ppwm/u_mem/_0245_ ),
    .C(\u_ppwm/u_mem/_0246_ ),
    .D(\u_ppwm/u_mem/_0248_ ),
    .Y(\u_ppwm/u_mem/_0249_ ));
 sg13g2_a21o_1 \u_ppwm/u_mem/_0738_  (.A2(\u_ppwm/u_mem/_0244_ ),
    .A1(net625),
    .B1(\u_ppwm/u_mem/_0249_ ),
    .X(\u_ppwm/u_mem/_0005_ ));
 sg13g2_nand3_1 \u_ppwm/u_mem/_0739_  (.B(net423),
    .C(net513),
    .A(net1),
    .Y(\u_ppwm/u_mem/_0250_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0740_  (.B1(\u_ppwm/u_mem/_0250_ ),
    .Y(\u_ppwm/u_mem/_0006_ ),
    .A1(net603),
    .A2(\u_ppwm/u_mem/_0248_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0741_  (.A0(\u_ppwm/u_mem/memory[70] ),
    .A1(\u_ppwm/u_mem/memory[77] ),
    .S(net411),
    .X(\u_ppwm/u_mem/_0251_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0742_  (.A0(\u_ppwm/u_mem/memory[56] ),
    .A1(\u_ppwm/u_mem/memory[63] ),
    .S(net413),
    .X(\u_ppwm/u_mem/_0252_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0743_  (.Y(\u_ppwm/u_mem/_0253_ ),
    .A(net334),
    .B(\u_ppwm/u_mem/_0252_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0744_  (.A1(net404),
    .A2(\u_ppwm/u_mem/_0251_ ),
    .Y(\u_ppwm/u_mem/_0254_ ),
    .B1(net403));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0745_  (.A0(\u_ppwm/u_mem/memory[84] ),
    .A1(\u_ppwm/u_mem/memory[91] ),
    .S(net410),
    .X(\u_ppwm/u_mem/_0255_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0746_  (.Y(\u_ppwm/u_mem/_0256_ ),
    .A(net334),
    .B(\u_ppwm/u_mem/_0255_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0747_  (.A0(\u_ppwm/u_mem/memory[98] ),
    .A1(\u_ppwm/u_mem/memory[105] ),
    .S(net410),
    .X(\u_ppwm/u_mem/_0257_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0748_  (.A1(net404),
    .A2(\u_ppwm/u_mem/_0257_ ),
    .Y(\u_ppwm/u_mem/_0258_ ),
    .B1(net333));
 sg13g2_a221oi_1 \u_ppwm/u_mem/_0749_  (.B2(\u_ppwm/u_mem/_0258_ ),
    .C1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0256_ ),
    .A1(\u_ppwm/u_mem/_0253_ ),
    .Y(\u_ppwm/u_mem/_0259_ ),
    .A2(\u_ppwm/u_mem/_0254_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0750_  (.S0(net417),
    .A0(\u_ppwm/u_mem/memory[0] ),
    .A1(\u_ppwm/u_mem/memory[7] ),
    .A2(\u_ppwm/u_mem/memory[14] ),
    .A3(\u_ppwm/u_mem/memory[21] ),
    .S1(net408),
    .X(\u_ppwm/u_mem/_0260_ ));
 sg13g2_nand2b_1 \u_ppwm/u_mem/_0751_  (.Y(\u_ppwm/u_mem/_0261_ ),
    .B(net332),
    .A_N(\u_ppwm/u_mem/_0260_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0752_  (.A0(\u_ppwm/u_mem/memory[42] ),
    .A1(\u_ppwm/u_mem/memory[49] ),
    .S(net416),
    .X(\u_ppwm/u_mem/_0262_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0753_  (.A0(\u_ppwm/u_mem/memory[28] ),
    .A1(\u_ppwm/u_mem/memory[35] ),
    .S(net415),
    .X(\u_ppwm/u_mem/_0263_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0754_  (.Y(\u_ppwm/u_mem/_0264_ ),
    .A(net335),
    .B(\u_ppwm/u_mem/_0263_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0755_  (.A1(net407),
    .A2(\u_ppwm/u_mem/_0262_ ),
    .Y(\u_ppwm/u_mem/_0265_ ),
    .B1(net332));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0756_  (.A1(\u_ppwm/u_mem/_0264_ ),
    .A2(\u_ppwm/u_mem/_0265_ ),
    .Y(\u_ppwm/u_mem/_0266_ ),
    .B1(net400));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0757_  (.A2(\u_ppwm/u_mem/_0266_ ),
    .A1(\u_ppwm/u_mem/_0261_ ),
    .B1(\u_ppwm/u_mem/_0259_ ),
    .X(\u_ppwm/instr[0] ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0758_  (.A0(\u_ppwm/u_mem/memory[99] ),
    .A1(\u_ppwm/u_mem/memory[106] ),
    .S(net410),
    .X(\u_ppwm/u_mem/_0267_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0759_  (.A0(\u_ppwm/u_mem/memory[85] ),
    .A1(\u_ppwm/u_mem/memory[92] ),
    .S(net412),
    .X(\u_ppwm/u_mem/_0268_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0760_  (.Y(\u_ppwm/u_mem/_0269_ ),
    .A(net334),
    .B(\u_ppwm/u_mem/_0268_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0761_  (.A1(net406),
    .A2(\u_ppwm/u_mem/_0267_ ),
    .Y(\u_ppwm/u_mem/_0270_ ),
    .B1(net333));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0762_  (.S0(net413),
    .A0(\u_ppwm/u_mem/memory[57] ),
    .A1(\u_ppwm/u_mem/memory[64] ),
    .A2(\u_ppwm/u_mem/memory[71] ),
    .A3(\u_ppwm/u_mem/memory[78] ),
    .S1(net406),
    .X(\u_ppwm/u_mem/_0271_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0763_  (.B1(net400),
    .Y(\u_ppwm/u_mem/_0272_ ),
    .A1(net403),
    .A2(\u_ppwm/u_mem/_0271_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0764_  (.A1(\u_ppwm/u_mem/_0269_ ),
    .A2(\u_ppwm/u_mem/_0270_ ),
    .Y(\u_ppwm/u_mem/_0273_ ),
    .B1(\u_ppwm/u_mem/_0272_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0765_  (.Y(\u_ppwm/u_mem/_0274_ ),
    .A(\u_ppwm/u_mem/memory[36] ),
    .B(net415));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0766_  (.B1(\u_ppwm/u_mem/_0274_ ),
    .Y(\u_ppwm/u_mem/_0275_ ),
    .A1(\u_ppwm/u_mem/_0209_ ),
    .A2(net417));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0767_  (.Y(\u_ppwm/u_mem/_0276_ ),
    .A(\u_ppwm/u_mem/memory[50] ),
    .B(net418));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0768_  (.B1(\u_ppwm/u_mem/_0276_ ),
    .Y(\u_ppwm/u_mem/_0277_ ),
    .A1(\u_ppwm/u_mem/_0195_ ),
    .A2(net418));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0769_  (.Y(\u_ppwm/u_mem/_0278_ ),
    .A(\u_ppwm/u_mem/memory[22] ),
    .B(net417));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0770_  (.B1(\u_ppwm/u_mem/_0278_ ),
    .Y(\u_ppwm/u_mem/_0279_ ),
    .A1(\u_ppwm/u_mem/_0223_ ),
    .A2(net417));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0771_  (.Y(\u_ppwm/u_mem/_0280_ ),
    .A(\u_ppwm/u_mem/memory[8] ),
    .B(net417));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0772_  (.B1(\u_ppwm/u_mem/_0280_ ),
    .Y(\u_ppwm/u_mem/_0281_ ),
    .A1(\u_ppwm/u_mem/_0237_ ),
    .A2(net420));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0773_  (.S0(net408),
    .A0(\u_ppwm/u_mem/_0275_ ),
    .A1(\u_ppwm/u_mem/_0277_ ),
    .A2(\u_ppwm/u_mem/_0281_ ),
    .A3(\u_ppwm/u_mem/_0279_ ),
    .S1(net332),
    .X(\u_ppwm/u_mem/_0282_ ));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0774_  (.A2(\u_ppwm/u_mem/_0282_ ),
    .A1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0273_ ),
    .X(\u_ppwm/instr[1] ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0775_  (.A0(\u_ppwm/u_mem/memory[100] ),
    .A1(\u_ppwm/u_mem/memory[107] ),
    .S(net410),
    .X(\u_ppwm/u_mem/_0283_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0776_  (.Y(\u_ppwm/u_mem/_0284_ ),
    .A(net404),
    .B(\u_ppwm/u_mem/_0283_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0777_  (.A0(\u_ppwm/u_mem/memory[86] ),
    .A1(\u_ppwm/u_mem/memory[93] ),
    .S(net413),
    .X(\u_ppwm/u_mem/_0285_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0778_  (.A1(net334),
    .A2(\u_ppwm/u_mem/_0285_ ),
    .Y(\u_ppwm/u_mem/_0286_ ),
    .B1(net333));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0779_  (.A0(\u_ppwm/u_mem/memory[72] ),
    .A1(\u_ppwm/u_mem/memory[79] ),
    .S(net411),
    .X(\u_ppwm/u_mem/_0287_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0780_  (.Y(\u_ppwm/u_mem/_0288_ ),
    .A(net405),
    .B(\u_ppwm/u_mem/_0287_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0781_  (.A0(\u_ppwm/u_mem/memory[58] ),
    .A1(\u_ppwm/u_mem/memory[65] ),
    .S(net411),
    .X(\u_ppwm/u_mem/_0289_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0782_  (.A1(net334),
    .A2(\u_ppwm/u_mem/_0289_ ),
    .Y(\u_ppwm/u_mem/_0290_ ),
    .B1(net403));
 sg13g2_a221oi_1 \u_ppwm/u_mem/_0783_  (.B2(\u_ppwm/u_mem/_0290_ ),
    .C1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0288_ ),
    .A1(\u_ppwm/u_mem/_0284_ ),
    .Y(\u_ppwm/u_mem/_0291_ ),
    .A2(\u_ppwm/u_mem/_0286_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0784_  (.Y(\u_ppwm/u_mem/_0292_ ),
    .A(\u_ppwm/u_mem/memory[37] ),
    .B(net418));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0785_  (.B1(\u_ppwm/u_mem/_0292_ ),
    .Y(\u_ppwm/u_mem/_0293_ ),
    .A1(\u_ppwm/u_mem/_0208_ ),
    .A2(net418));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0786_  (.Y(\u_ppwm/u_mem/_0294_ ),
    .A(\u_ppwm/u_mem/memory[51] ),
    .B(net419));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0787_  (.B1(\u_ppwm/u_mem/_0294_ ),
    .Y(\u_ppwm/u_mem/_0295_ ),
    .A1(\u_ppwm/u_mem/_0194_ ),
    .A2(net419));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0788_  (.Y(\u_ppwm/u_mem/_0296_ ),
    .A(\u_ppwm/u_mem/memory[23] ),
    .B(net419));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0789_  (.B1(\u_ppwm/u_mem/_0296_ ),
    .Y(\u_ppwm/u_mem/_0297_ ),
    .A1(\u_ppwm/u_mem/_0222_ ),
    .A2(net418));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0790_  (.Y(\u_ppwm/u_mem/_0298_ ),
    .A(\u_ppwm/u_mem/memory[9] ),
    .B(net417));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0791_  (.B1(\u_ppwm/u_mem/_0298_ ),
    .Y(\u_ppwm/u_mem/_0299_ ),
    .A1(\u_ppwm/u_mem/_0236_ ),
    .A2(net418));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0792_  (.S0(net408),
    .A0(\u_ppwm/u_mem/_0293_ ),
    .A1(\u_ppwm/u_mem/_0295_ ),
    .A2(\u_ppwm/u_mem/_0299_ ),
    .A3(\u_ppwm/u_mem/_0297_ ),
    .S1(\u_ppwm/u_mem/_0241_ ),
    .X(\u_ppwm/u_mem/_0300_ ));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0793_  (.A2(\u_ppwm/u_mem/_0300_ ),
    .A1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0291_ ),
    .X(\u_ppwm/instr[2] ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0794_  (.A0(\u_ppwm/u_mem/memory[101] ),
    .A1(\u_ppwm/u_mem/_0000_ ),
    .S(net410),
    .X(\u_ppwm/u_mem/_0301_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0795_  (.Y(\u_ppwm/u_mem/_0302_ ),
    .A(net404),
    .B(\u_ppwm/u_mem/_0301_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0796_  (.A0(\u_ppwm/u_mem/memory[87] ),
    .A1(\u_ppwm/u_mem/memory[94] ),
    .S(net413),
    .X(\u_ppwm/u_mem/_0303_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0797_  (.A1(net334),
    .A2(\u_ppwm/u_mem/_0303_ ),
    .Y(\u_ppwm/u_mem/_0304_ ),
    .B1(net333));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0798_  (.A0(\u_ppwm/u_mem/memory[73] ),
    .A1(\u_ppwm/u_mem/memory[80] ),
    .S(net414),
    .X(\u_ppwm/u_mem/_0305_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0799_  (.Y(\u_ppwm/u_mem/_0306_ ),
    .A(net405),
    .B(\u_ppwm/u_mem/_0305_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0800_  (.A0(\u_ppwm/u_mem/memory[59] ),
    .A1(\u_ppwm/u_mem/memory[66] ),
    .S(net411),
    .X(\u_ppwm/u_mem/_0307_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0801_  (.A1(net335),
    .A2(\u_ppwm/u_mem/_0307_ ),
    .Y(\u_ppwm/u_mem/_0308_ ),
    .B1(net403));
 sg13g2_a221oi_1 \u_ppwm/u_mem/_0802_  (.B2(\u_ppwm/u_mem/_0308_ ),
    .C1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0306_ ),
    .A1(\u_ppwm/u_mem/_0302_ ),
    .Y(\u_ppwm/u_mem/_0309_ ),
    .A2(\u_ppwm/u_mem/_0304_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0803_  (.A0(\u_ppwm/u_mem/_0207_ ),
    .A1(\u_ppwm/u_mem/_0200_ ),
    .S(net416),
    .X(\u_ppwm/u_mem/_0310_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0804_  (.A0(\u_ppwm/u_mem/memory[45] ),
    .A1(\u_ppwm/u_mem/memory[52] ),
    .S(net418),
    .X(\u_ppwm/u_mem/_0311_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0805_  (.A1(net409),
    .A2(\u_ppwm/u_mem/_0311_ ),
    .Y(\u_ppwm/u_mem/_0312_ ),
    .B1(net332));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0806_  (.B1(\u_ppwm/u_mem/_0312_ ),
    .Y(\u_ppwm/u_mem/_0313_ ),
    .A1(net407),
    .A2(\u_ppwm/u_mem/_0310_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0807_  (.S0(net335),
    .A0(\u_ppwm/u_mem/_0221_ ),
    .A1(\u_ppwm/u_mem/_0235_ ),
    .A2(\u_ppwm/u_mem/_0214_ ),
    .A3(\u_ppwm/u_mem/_0228_ ),
    .S1(net419),
    .X(\u_ppwm/u_mem/_0314_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0808_  (.A1(net332),
    .A2(\u_ppwm/u_mem/_0314_ ),
    .Y(\u_ppwm/u_mem/_0315_ ),
    .B1(net401));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0809_  (.A2(\u_ppwm/u_mem/_0315_ ),
    .A1(\u_ppwm/u_mem/_0313_ ),
    .B1(\u_ppwm/u_mem/_0309_ ),
    .X(\u_ppwm/instr[3] ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0810_  (.B1(net404),
    .Y(\u_ppwm/u_mem/_0316_ ),
    .A1(\u_ppwm/u_mem/memory[102] ),
    .A2(net411));
 sg13g2_a21o_1 \u_ppwm/u_mem/_0811_  (.A2(net412),
    .A1(\u_ppwm/u_mem/_0129_ ),
    .B1(\u_ppwm/u_mem/_0316_ ),
    .X(\u_ppwm/u_mem/_0317_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0812_  (.A0(\u_ppwm/u_mem/memory[88] ),
    .A1(\u_ppwm/u_mem/memory[95] ),
    .S(net412),
    .X(\u_ppwm/u_mem/_0318_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0813_  (.A1(net334),
    .A2(\u_ppwm/u_mem/_0318_ ),
    .Y(\u_ppwm/u_mem/_0319_ ),
    .B1(net333));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0814_  (.S0(net411),
    .A0(\u_ppwm/u_mem/memory[60] ),
    .A1(\u_ppwm/u_mem/memory[67] ),
    .A2(\u_ppwm/u_mem/memory[74] ),
    .A3(\u_ppwm/u_mem/memory[81] ),
    .S1(net405),
    .X(\u_ppwm/u_mem/_0320_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0815_  (.B1(net400),
    .Y(\u_ppwm/u_mem/_0321_ ),
    .A1(net403),
    .A2(\u_ppwm/u_mem/_0320_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0816_  (.A1(\u_ppwm/u_mem/_0317_ ),
    .A2(\u_ppwm/u_mem/_0319_ ),
    .Y(\u_ppwm/u_mem/_0322_ ),
    .B1(\u_ppwm/u_mem/_0321_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0817_  (.A0(\u_ppwm/u_mem/memory[18] ),
    .A1(\u_ppwm/u_mem/memory[25] ),
    .S(net418),
    .X(\u_ppwm/u_mem/_0323_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0818_  (.Y(\u_ppwm/u_mem/_0324_ ),
    .A(net409),
    .B(\u_ppwm/u_mem/_0323_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0819_  (.A0(\u_ppwm/u_mem/memory[4] ),
    .A1(\u_ppwm/u_mem/memory[11] ),
    .S(net417),
    .X(\u_ppwm/u_mem/_0325_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0820_  (.A1(net335),
    .A2(\u_ppwm/u_mem/_0325_ ),
    .Y(\u_ppwm/u_mem/_0326_ ),
    .B1(\u_ppwm/pc[2] ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0821_  (.B1(net408),
    .Y(\u_ppwm/u_mem/_0327_ ),
    .A1(\u_ppwm/u_mem/memory[46] ),
    .A2(net415));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0822_  (.A1(\u_ppwm/u_mem/_0185_ ),
    .A2(net416),
    .Y(\u_ppwm/u_mem/_0328_ ),
    .B1(\u_ppwm/u_mem/_0327_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0823_  (.A0(\u_ppwm/u_mem/memory[32] ),
    .A1(\u_ppwm/u_mem/memory[39] ),
    .S(net416),
    .X(\u_ppwm/u_mem/_0329_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0824_  (.A1(net335),
    .A2(\u_ppwm/u_mem/_0329_ ),
    .Y(\u_ppwm/u_mem/_0330_ ),
    .B1(net332));
 sg13g2_nand2b_1 \u_ppwm/u_mem/_0825_  (.Y(\u_ppwm/u_mem/_0331_ ),
    .B(\u_ppwm/u_mem/_0330_ ),
    .A_N(\u_ppwm/u_mem/_0328_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0826_  (.A1(\u_ppwm/u_mem/_0324_ ),
    .A2(\u_ppwm/u_mem/_0326_ ),
    .Y(\u_ppwm/u_mem/_0332_ ),
    .B1(net401));
 sg13g2_a21o_1 \u_ppwm/u_mem/_0827_  (.A2(\u_ppwm/u_mem/_0332_ ),
    .A1(\u_ppwm/u_mem/_0331_ ),
    .B1(\u_ppwm/u_mem/_0322_ ),
    .X(\u_ppwm/instr[4] ));
 sg13g2_nor2b_1 \u_ppwm/u_mem/_0828_  (.A(\u_ppwm/u_mem/_0002_ ),
    .B_N(net412),
    .Y(\u_ppwm/u_mem/_0333_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0829_  (.B1(net404),
    .Y(\u_ppwm/u_mem/_0334_ ),
    .A1(\u_ppwm/u_mem/memory[103] ),
    .A2(net412));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0830_  (.Y(\u_ppwm/u_mem/_0335_ ),
    .A(\u_ppwm/u_mem/memory[96] ),
    .B(net412));
 sg13g2_nand2b_1 \u_ppwm/u_mem/_0831_  (.Y(\u_ppwm/u_mem/_0336_ ),
    .B(\u_ppwm/u_mem/memory[89] ),
    .A_N(net412));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0832_  (.A1(\u_ppwm/u_mem/_0335_ ),
    .A2(\u_ppwm/u_mem/_0336_ ),
    .Y(\u_ppwm/u_mem/_0337_ ),
    .B1(net406));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0833_  (.B1(net403),
    .Y(\u_ppwm/u_mem/_0338_ ),
    .A1(\u_ppwm/u_mem/_0333_ ),
    .A2(\u_ppwm/u_mem/_0334_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0834_  (.S0(net414),
    .A0(\u_ppwm/u_mem/memory[61] ),
    .A1(\u_ppwm/u_mem/memory[68] ),
    .A2(\u_ppwm/u_mem/memory[75] ),
    .A3(\u_ppwm/u_mem/memory[82] ),
    .S1(net405),
    .X(\u_ppwm/u_mem/_0339_ ));
 sg13g2_nor2_1 \u_ppwm/u_mem/_0835_  (.A(net403),
    .B(\u_ppwm/u_mem/_0339_ ),
    .Y(\u_ppwm/u_mem/_0340_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0836_  (.B1(net400),
    .Y(\u_ppwm/u_mem/_0341_ ),
    .A1(\u_ppwm/u_mem/_0337_ ),
    .A2(\u_ppwm/u_mem/_0338_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0837_  (.A0(\u_ppwm/u_mem/memory[33] ),
    .A1(\u_ppwm/u_mem/memory[40] ),
    .S(net416),
    .X(\u_ppwm/u_mem/_0342_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0838_  (.A0(\u_ppwm/u_mem/memory[47] ),
    .A1(\u_ppwm/u_mem/memory[54] ),
    .S(net416),
    .X(\u_ppwm/u_mem/_0343_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0839_  (.A0(\u_ppwm/u_mem/memory[19] ),
    .A1(\u_ppwm/u_mem/memory[26] ),
    .S(net415),
    .X(\u_ppwm/u_mem/_0344_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0840_  (.A0(\u_ppwm/u_mem/memory[5] ),
    .A1(\u_ppwm/u_mem/memory[12] ),
    .S(net415),
    .X(\u_ppwm/u_mem/_0345_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0841_  (.S0(net407),
    .A0(\u_ppwm/u_mem/_0342_ ),
    .A1(\u_ppwm/u_mem/_0343_ ),
    .A2(\u_ppwm/u_mem/_0345_ ),
    .A3(\u_ppwm/u_mem/_0344_ ),
    .S1(net332),
    .X(\u_ppwm/u_mem/_0346_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0842_  (.Y(\u_ppwm/u_mem/_0347_ ),
    .A(\u_ppwm/u_mem/_0242_ ),
    .B(\u_ppwm/u_mem/_0346_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0843_  (.B1(\u_ppwm/u_mem/_0347_ ),
    .Y(\u_ppwm/instr[5] ),
    .A1(\u_ppwm/u_mem/_0340_ ),
    .A2(\u_ppwm/u_mem/_0341_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0844_  (.A0(\u_ppwm/u_mem/memory[76] ),
    .A1(\u_ppwm/u_mem/memory[83] ),
    .S(net410),
    .X(\u_ppwm/u_mem/_0348_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0845_  (.Y(\u_ppwm/u_mem/_0349_ ),
    .A(net404),
    .B(\u_ppwm/u_mem/_0348_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0846_  (.A0(\u_ppwm/u_mem/memory[62] ),
    .A1(\u_ppwm/u_mem/memory[69] ),
    .S(net411),
    .X(\u_ppwm/u_mem/_0350_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0847_  (.A1(net335),
    .A2(\u_ppwm/u_mem/_0350_ ),
    .Y(\u_ppwm/u_mem/_0351_ ),
    .B1(net403));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0848_  (.A0(\u_ppwm/u_mem/memory[90] ),
    .A1(\u_ppwm/u_mem/memory[97] ),
    .S(net410),
    .X(\u_ppwm/u_mem/_0352_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0849_  (.A0(\u_ppwm/u_mem/memory[104] ),
    .A1(\u_ppwm/u_mem/_0003_ ),
    .S(net410),
    .X(\u_ppwm/u_mem/_0353_ ));
 sg13g2_nand2_1 \u_ppwm/u_mem/_0850_  (.Y(\u_ppwm/u_mem/_0354_ ),
    .A(net404),
    .B(\u_ppwm/u_mem/_0353_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0851_  (.A1(net334),
    .A2(\u_ppwm/u_mem/_0352_ ),
    .Y(\u_ppwm/u_mem/_0355_ ),
    .B1(net333));
 sg13g2_a221oi_1 \u_ppwm/u_mem/_0852_  (.B2(\u_ppwm/u_mem/_0355_ ),
    .C1(\u_ppwm/u_mem/_0242_ ),
    .B1(\u_ppwm/u_mem/_0354_ ),
    .A1(\u_ppwm/u_mem/_0349_ ),
    .Y(\u_ppwm/u_mem/_0356_ ),
    .A2(\u_ppwm/u_mem/_0351_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0853_  (.A0(\u_ppwm/u_mem/_0204_ ),
    .A1(\u_ppwm/u_mem/_0197_ ),
    .S(net416),
    .X(\u_ppwm/u_mem/_0357_ ));
 sg13g2_mux2_1 \u_ppwm/u_mem/_0854_  (.A0(\u_ppwm/u_mem/memory[48] ),
    .A1(\u_ppwm/u_mem/memory[55] ),
    .S(net413),
    .X(\u_ppwm/u_mem/_0358_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0855_  (.A1(net408),
    .A2(\u_ppwm/u_mem/_0358_ ),
    .Y(\u_ppwm/u_mem/_0359_ ),
    .B1(net333));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0856_  (.B1(\u_ppwm/u_mem/_0359_ ),
    .Y(\u_ppwm/u_mem/_0360_ ),
    .A1(net408),
    .A2(\u_ppwm/u_mem/_0357_ ));
 sg13g2_mux4_1 \u_ppwm/u_mem/_0857_  (.S0(net335),
    .A0(\u_ppwm/u_mem/_0218_ ),
    .A1(\u_ppwm/u_mem/_0232_ ),
    .A2(\u_ppwm/u_mem/_0211_ ),
    .A3(\u_ppwm/u_mem/_0225_ ),
    .S1(net417),
    .X(\u_ppwm/u_mem/_0361_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0858_  (.A1(net332),
    .A2(\u_ppwm/u_mem/_0361_ ),
    .Y(\u_ppwm/u_mem/_0362_ ),
    .B1(net401));
 sg13g2_a21o_2 \u_ppwm/u_mem/_0859_  (.A2(\u_ppwm/u_mem/_0362_ ),
    .A1(\u_ppwm/u_mem/_0360_ ),
    .B1(\u_ppwm/u_mem/_0356_ ),
    .X(\u_ppwm/instr[6] ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0860_  (.B1(net447),
    .Y(\u_ppwm/u_mem/_0363_ ),
    .A1(net360),
    .A2(\u_ppwm/u_mem/memory[0] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0861_  (.A1(net360),
    .A2(\u_ppwm/u_mem/_0237_ ),
    .Y(\u_ppwm/u_mem/_0007_ ),
    .B1(\u_ppwm/u_mem/_0363_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0862_  (.B1(net451),
    .Y(\u_ppwm/u_mem/_0364_ ),
    .A1(net361),
    .A2(net511));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0863_  (.A1(net361),
    .A2(\u_ppwm/u_mem/_0236_ ),
    .Y(\u_ppwm/u_mem/_0008_ ),
    .B1(\u_ppwm/u_mem/_0364_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0864_  (.B1(net450),
    .Y(\u_ppwm/u_mem/_0365_ ),
    .A1(net370),
    .A2(\u_ppwm/u_mem/memory[2] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0865_  (.A1(net370),
    .A2(\u_ppwm/u_mem/_0235_ ),
    .Y(\u_ppwm/u_mem/_0009_ ),
    .B1(\u_ppwm/u_mem/_0365_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0866_  (.B1(net450),
    .Y(\u_ppwm/u_mem/_0366_ ),
    .A1(net370),
    .A2(net501));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0867_  (.A1(net370),
    .A2(\u_ppwm/u_mem/_0234_ ),
    .Y(\u_ppwm/u_mem/_0010_ ),
    .B1(\u_ppwm/u_mem/_0366_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0868_  (.B1(net448),
    .Y(\u_ppwm/u_mem/_0367_ ),
    .A1(net362),
    .A2(net527));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0869_  (.A1(net362),
    .A2(\u_ppwm/u_mem/_0233_ ),
    .Y(\u_ppwm/u_mem/_0011_ ),
    .B1(\u_ppwm/u_mem/_0367_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0870_  (.B1(net443),
    .Y(\u_ppwm/u_mem/_0368_ ),
    .A1(net358),
    .A2(net532));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0871_  (.A1(net359),
    .A2(\u_ppwm/u_mem/_0232_ ),
    .Y(\u_ppwm/u_mem/_0012_ ),
    .B1(\u_ppwm/u_mem/_0368_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0872_  (.B1(net448),
    .Y(\u_ppwm/u_mem/_0369_ ),
    .A1(net363),
    .A2(\u_ppwm/u_mem/memory[6] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0873_  (.A1(net363),
    .A2(\u_ppwm/u_mem/_0231_ ),
    .Y(\u_ppwm/u_mem/_0013_ ),
    .B1(\u_ppwm/u_mem/_0369_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0874_  (.B1(net447),
    .Y(\u_ppwm/u_mem/_0370_ ),
    .A1(net363),
    .A2(net481));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0875_  (.A1(net360),
    .A2(\u_ppwm/u_mem/_0230_ ),
    .Y(\u_ppwm/u_mem/_0014_ ),
    .B1(\u_ppwm/u_mem/_0370_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0876_  (.B1(net447),
    .Y(\u_ppwm/u_mem/_0371_ ),
    .A1(net360),
    .A2(\u_ppwm/u_mem/memory[8] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0877_  (.A1(net361),
    .A2(\u_ppwm/u_mem/_0229_ ),
    .Y(\u_ppwm/u_mem/_0015_ ),
    .B1(\u_ppwm/u_mem/_0371_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0878_  (.B1(net447),
    .Y(\u_ppwm/u_mem/_0372_ ),
    .A1(net371),
    .A2(net241));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0879_  (.A1(net370),
    .A2(\u_ppwm/u_mem/_0228_ ),
    .Y(\u_ppwm/u_mem/_0016_ ),
    .B1(\u_ppwm/u_mem/_0372_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0880_  (.B1(net447),
    .Y(\u_ppwm/u_mem/_0373_ ),
    .A1(net371),
    .A2(\u_ppwm/u_mem/memory[10] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0881_  (.A1(net370),
    .A2(\u_ppwm/u_mem/_0227_ ),
    .Y(\u_ppwm/u_mem/_0017_ ),
    .B1(\u_ppwm/u_mem/_0373_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0882_  (.B1(net448),
    .Y(\u_ppwm/u_mem/_0374_ ),
    .A1(net362),
    .A2(net464));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0883_  (.A1(net362),
    .A2(\u_ppwm/u_mem/_0226_ ),
    .Y(\u_ppwm/u_mem/_0018_ ),
    .B1(\u_ppwm/u_mem/_0374_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0884_  (.B1(net448),
    .Y(\u_ppwm/u_mem/_0375_ ),
    .A1(net359),
    .A2(net469));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0885_  (.A1(net359),
    .A2(\u_ppwm/u_mem/_0225_ ),
    .Y(\u_ppwm/u_mem/_0019_ ),
    .B1(\u_ppwm/u_mem/_0375_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0886_  (.B1(net448),
    .Y(\u_ppwm/u_mem/_0376_ ),
    .A1(net362),
    .A2(net491));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0887_  (.A1(net362),
    .A2(\u_ppwm/u_mem/_0224_ ),
    .Y(\u_ppwm/u_mem/_0020_ ),
    .B1(\u_ppwm/u_mem/_0376_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0888_  (.B1(net447),
    .Y(\u_ppwm/u_mem/_0377_ ),
    .A1(net360),
    .A2(net506));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0889_  (.A1(net360),
    .A2(\u_ppwm/u_mem/_0223_ ),
    .Y(\u_ppwm/u_mem/_0021_ ),
    .B1(\u_ppwm/u_mem/_0377_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0890_  (.B1(net447),
    .Y(\u_ppwm/u_mem/_0378_ ),
    .A1(net370),
    .A2(net589));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0891_  (.A1(net370),
    .A2(\u_ppwm/u_mem/_0222_ ),
    .Y(\u_ppwm/u_mem/_0022_ ),
    .B1(\u_ppwm/u_mem/_0378_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0892_  (.B1(net450),
    .Y(\u_ppwm/u_mem/_0379_ ),
    .A1(net371),
    .A2(\u_ppwm/u_mem/memory[16] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0893_  (.A1(net372),
    .A2(\u_ppwm/u_mem/_0221_ ),
    .Y(\u_ppwm/u_mem/_0023_ ),
    .B1(\u_ppwm/u_mem/_0379_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0894_  (.B1(net450),
    .Y(\u_ppwm/u_mem/_0380_ ),
    .A1(net371),
    .A2(\u_ppwm/u_mem/memory[17] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0895_  (.A1(net371),
    .A2(\u_ppwm/u_mem/_0220_ ),
    .Y(\u_ppwm/u_mem/_0024_ ),
    .B1(\u_ppwm/u_mem/_0380_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0896_  (.B1(net449),
    .Y(\u_ppwm/u_mem/_0381_ ),
    .A1(net372),
    .A2(net301));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0897_  (.A1(net372),
    .A2(\u_ppwm/u_mem/_0219_ ),
    .Y(\u_ppwm/u_mem/_0025_ ),
    .B1(\u_ppwm/u_mem/_0381_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0898_  (.B1(net443),
    .Y(\u_ppwm/u_mem/_0382_ ),
    .A1(net358),
    .A2(net503));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0899_  (.A1(net358),
    .A2(\u_ppwm/u_mem/_0218_ ),
    .Y(\u_ppwm/u_mem/_0026_ ),
    .B1(\u_ppwm/u_mem/_0382_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0900_  (.B1(net448),
    .Y(\u_ppwm/u_mem/_0383_ ),
    .A1(net362),
    .A2(\u_ppwm/u_mem/memory[20] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0901_  (.A1(net362),
    .A2(\u_ppwm/u_mem/_0217_ ),
    .Y(\u_ppwm/u_mem/_0027_ ),
    .B1(\u_ppwm/u_mem/_0383_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0902_  (.B1(net447),
    .Y(\u_ppwm/u_mem/_0384_ ),
    .A1(net360),
    .A2(net479));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0903_  (.A1(net360),
    .A2(\u_ppwm/u_mem/_0216_ ),
    .Y(\u_ppwm/u_mem/_0028_ ),
    .B1(\u_ppwm/u_mem/_0384_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0904_  (.B1(net448),
    .Y(\u_ppwm/u_mem/_0385_ ),
    .A1(net361),
    .A2(net500));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0905_  (.A1(net361),
    .A2(\u_ppwm/u_mem/_0215_ ),
    .Y(\u_ppwm/u_mem/_0029_ ),
    .B1(\u_ppwm/u_mem/_0385_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0906_  (.B1(net450),
    .Y(\u_ppwm/u_mem/_0386_ ),
    .A1(net372),
    .A2(\u_ppwm/u_mem/memory[23] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0907_  (.A1(net372),
    .A2(\u_ppwm/u_mem/_0214_ ),
    .Y(\u_ppwm/u_mem/_0030_ ),
    .B1(\u_ppwm/u_mem/_0386_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0908_  (.B1(net450),
    .Y(\u_ppwm/u_mem/_0387_ ),
    .A1(net371),
    .A2(\u_ppwm/u_mem/memory[24] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0909_  (.A1(net371),
    .A2(\u_ppwm/u_mem/_0213_ ),
    .Y(\u_ppwm/u_mem/_0031_ ),
    .B1(\u_ppwm/u_mem/_0387_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0910_  (.B1(net449),
    .Y(\u_ppwm/u_mem/_0388_ ),
    .A1(net372),
    .A2(net299));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0911_  (.A1(net372),
    .A2(\u_ppwm/u_mem/_0212_ ),
    .Y(\u_ppwm/u_mem/_0032_ ),
    .B1(\u_ppwm/u_mem/_0388_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0912_  (.B1(net443),
    .Y(\u_ppwm/u_mem/_0389_ ),
    .A1(net358),
    .A2(\u_ppwm/u_mem/memory[26] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0913_  (.A1(net359),
    .A2(\u_ppwm/u_mem/_0211_ ),
    .Y(\u_ppwm/u_mem/_0033_ ),
    .B1(\u_ppwm/u_mem/_0389_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0914_  (.B1(net446),
    .Y(\u_ppwm/u_mem/_0390_ ),
    .A1(net358),
    .A2(\u_ppwm/u_mem/memory[27] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0915_  (.A1(net358),
    .A2(\u_ppwm/u_mem/_0210_ ),
    .Y(\u_ppwm/u_mem/_0034_ ),
    .B1(\u_ppwm/u_mem/_0390_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0916_  (.B1(net446),
    .Y(\u_ppwm/u_mem/_0391_ ),
    .A1(net358),
    .A2(net235));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0917_  (.A1(net358),
    .A2(\u_ppwm/u_mem/_0209_ ),
    .Y(\u_ppwm/u_mem/_0035_ ),
    .B1(\u_ppwm/u_mem/_0391_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0918_  (.B1(net449),
    .Y(\u_ppwm/u_mem/_0392_ ),
    .A1(net365),
    .A2(\u_ppwm/u_mem/memory[29] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0919_  (.A1(net365),
    .A2(\u_ppwm/u_mem/_0208_ ),
    .Y(\u_ppwm/u_mem/_0036_ ),
    .B1(\u_ppwm/u_mem/_0392_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0920_  (.B1(net445),
    .Y(\u_ppwm/u_mem/_0393_ ),
    .A1(net368),
    .A2(\u_ppwm/u_mem/memory[30] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0921_  (.A1(net368),
    .A2(\u_ppwm/u_mem/_0207_ ),
    .Y(\u_ppwm/u_mem/_0037_ ),
    .B1(\u_ppwm/u_mem/_0393_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0922_  (.B1(net444),
    .Y(\u_ppwm/u_mem/_0394_ ),
    .A1(net366),
    .A2(\u_ppwm/u_mem/memory[31] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0923_  (.A1(net366),
    .A2(\u_ppwm/u_mem/_0206_ ),
    .Y(\u_ppwm/u_mem/_0038_ ),
    .B1(\u_ppwm/u_mem/_0394_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0924_  (.B1(net445),
    .Y(\u_ppwm/u_mem/_0395_ ),
    .A1(net366),
    .A2(net216));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0925_  (.A1(net356),
    .A2(\u_ppwm/u_mem/_0205_ ),
    .Y(\u_ppwm/u_mem/_0039_ ),
    .B1(\u_ppwm/u_mem/_0395_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0926_  (.B1(net444),
    .Y(\u_ppwm/u_mem/_0396_ ),
    .A1(net364),
    .A2(net272));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0927_  (.A1(net364),
    .A2(\u_ppwm/u_mem/_0204_ ),
    .Y(\u_ppwm/u_mem/_0040_ ),
    .B1(\u_ppwm/u_mem/_0396_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0928_  (.B1(net444),
    .Y(\u_ppwm/u_mem/_0397_ ),
    .A1(net364),
    .A2(\u_ppwm/u_mem/memory[34] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0929_  (.A1(net364),
    .A2(\u_ppwm/u_mem/_0203_ ),
    .Y(\u_ppwm/u_mem/_0041_ ),
    .B1(\u_ppwm/u_mem/_0397_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0930_  (.B1(net443),
    .Y(\u_ppwm/u_mem/_0398_ ),
    .A1(net364),
    .A2(net289));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0931_  (.A1(net364),
    .A2(\u_ppwm/u_mem/_0202_ ),
    .Y(\u_ppwm/u_mem/_0042_ ),
    .B1(\u_ppwm/u_mem/_0398_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0932_  (.B1(net445),
    .Y(\u_ppwm/u_mem/_0399_ ),
    .A1(net365),
    .A2(\u_ppwm/u_mem/memory[36] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0933_  (.A1(net365),
    .A2(\u_ppwm/u_mem/_0201_ ),
    .Y(\u_ppwm/u_mem/_0043_ ),
    .B1(\u_ppwm/u_mem/_0399_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0934_  (.B1(net445),
    .Y(\u_ppwm/u_mem/_0400_ ),
    .A1(net365),
    .A2(net459));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0935_  (.A1(net365),
    .A2(\u_ppwm/u_mem/_0200_ ),
    .Y(\u_ppwm/u_mem/_0044_ ),
    .B1(\u_ppwm/u_mem/_0400_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0936_  (.B1(net446),
    .Y(\u_ppwm/u_mem/_0401_ ),
    .A1(net366),
    .A2(\u_ppwm/u_mem/memory[38] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0937_  (.A1(net366),
    .A2(\u_ppwm/u_mem/_0199_ ),
    .Y(\u_ppwm/u_mem/_0045_ ),
    .B1(\u_ppwm/u_mem/_0401_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0938_  (.B1(net444),
    .Y(\u_ppwm/u_mem/_0402_ ),
    .A1(net366),
    .A2(net280));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0939_  (.A1(net366),
    .A2(\u_ppwm/u_mem/_0198_ ),
    .Y(\u_ppwm/u_mem/_0046_ ),
    .B1(\u_ppwm/u_mem/_0402_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0940_  (.B1(net444),
    .Y(\u_ppwm/u_mem/_0403_ ),
    .A1(net364),
    .A2(\u_ppwm/u_mem/memory[40] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0941_  (.A1(net364),
    .A2(\u_ppwm/u_mem/_0197_ ),
    .Y(\u_ppwm/u_mem/_0047_ ),
    .B1(\u_ppwm/u_mem/_0403_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0942_  (.B1(net445),
    .Y(\u_ppwm/u_mem/_0404_ ),
    .A1(net368),
    .A2(\u_ppwm/u_mem/memory[41] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0943_  (.A1(net368),
    .A2(\u_ppwm/u_mem/_0196_ ),
    .Y(\u_ppwm/u_mem/_0048_ ),
    .B1(\u_ppwm/u_mem/_0404_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0944_  (.B1(net449),
    .Y(\u_ppwm/u_mem/_0405_ ),
    .A1(net373),
    .A2(\u_ppwm/u_mem/memory[42] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0945_  (.A1(net373),
    .A2(\u_ppwm/u_mem/_0195_ ),
    .Y(\u_ppwm/u_mem/_0049_ ),
    .B1(\u_ppwm/u_mem/_0405_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0946_  (.B1(net450),
    .Y(\u_ppwm/u_mem/_0406_ ),
    .A1(net374),
    .A2(net519));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0947_  (.A1(net374),
    .A2(\u_ppwm/u_mem/_0194_ ),
    .Y(\u_ppwm/u_mem/_0050_ ),
    .B1(\u_ppwm/u_mem/_0406_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0948_  (.B1(net450),
    .Y(\u_ppwm/u_mem/_0407_ ),
    .A1(net373),
    .A2(\u_ppwm/u_mem/memory[44] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0949_  (.A1(net373),
    .A2(\u_ppwm/u_mem/_0193_ ),
    .Y(\u_ppwm/u_mem/_0051_ ),
    .B1(\u_ppwm/u_mem/_0407_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0950_  (.B1(net449),
    .Y(\u_ppwm/u_mem/_0408_ ),
    .A1(net374),
    .A2(net297));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0951_  (.A1(net368),
    .A2(\u_ppwm/u_mem/_0192_ ),
    .Y(\u_ppwm/u_mem/_0052_ ),
    .B1(\u_ppwm/u_mem/_0408_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0952_  (.B1(net445),
    .Y(\u_ppwm/u_mem/_0409_ ),
    .A1(net369),
    .A2(\u_ppwm/u_mem/memory[46] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0953_  (.A1(net369),
    .A2(\u_ppwm/u_mem/_0191_ ),
    .Y(\u_ppwm/u_mem/_0053_ ),
    .B1(\u_ppwm/u_mem/_0409_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0954_  (.B1(net444),
    .Y(\u_ppwm/u_mem/_0410_ ),
    .A1(net366),
    .A2(\u_ppwm/u_mem/memory[47] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0955_  (.A1(net367),
    .A2(\u_ppwm/u_mem/_0190_ ),
    .Y(\u_ppwm/u_mem/_0054_ ),
    .B1(\u_ppwm/u_mem/_0410_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0956_  (.B1(net444),
    .Y(\u_ppwm/u_mem/_0411_ ),
    .A1(net367),
    .A2(net247));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0957_  (.A1(net367),
    .A2(\u_ppwm/u_mem/_0189_ ),
    .Y(\u_ppwm/u_mem/_0055_ ),
    .B1(\u_ppwm/u_mem/_0411_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0958_  (.B1(net449),
    .Y(\u_ppwm/u_mem/_0412_ ),
    .A1(net368),
    .A2(\u_ppwm/u_mem/memory[49] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0959_  (.A1(net373),
    .A2(\u_ppwm/u_mem/_0188_ ),
    .Y(\u_ppwm/u_mem/_0056_ ),
    .B1(\u_ppwm/u_mem/_0412_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0960_  (.B1(net449),
    .Y(\u_ppwm/u_mem/_0413_ ),
    .A1(net373),
    .A2(\u_ppwm/u_mem/memory[50] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0961_  (.A1(net373),
    .A2(\u_ppwm/u_mem/_0187_ ),
    .Y(\u_ppwm/u_mem/_0057_ ),
    .B1(\u_ppwm/u_mem/_0413_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0962_  (.B1(net449),
    .Y(\u_ppwm/u_mem/_0414_ ),
    .A1(net373),
    .A2(net237));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0963_  (.A1(net374),
    .A2(\u_ppwm/u_mem/_0186_ ),
    .Y(\u_ppwm/u_mem/_0058_ ),
    .B1(\u_ppwm/u_mem/_0414_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0964_  (.B1(net445),
    .Y(\u_ppwm/u_mem/_0415_ ),
    .A1(net368),
    .A2(net306));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0965_  (.A1(net368),
    .A2(\u_ppwm/u_mem/_0185_ ),
    .Y(\u_ppwm/u_mem/_0059_ ),
    .B1(\u_ppwm/u_mem/_0415_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0966_  (.B1(net446),
    .Y(\u_ppwm/u_mem/_0416_ ),
    .A1(net369),
    .A2(\u_ppwm/u_mem/memory[53] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0967_  (.A1(net367),
    .A2(\u_ppwm/u_mem/_0184_ ),
    .Y(\u_ppwm/u_mem/_0060_ ),
    .B1(\u_ppwm/u_mem/_0416_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0968_  (.B1(net444),
    .Y(\u_ppwm/u_mem/_0417_ ),
    .A1(net367),
    .A2(net256));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0969_  (.A1(net367),
    .A2(\u_ppwm/u_mem/_0183_ ),
    .Y(\u_ppwm/u_mem/_0061_ ),
    .B1(\u_ppwm/u_mem/_0417_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0970_  (.B1(net435),
    .Y(\u_ppwm/u_mem/_0418_ ),
    .A1(net356),
    .A2(\u_ppwm/u_mem/memory[55] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0971_  (.A1(net356),
    .A2(\u_ppwm/u_mem/_0182_ ),
    .Y(\u_ppwm/u_mem/_0062_ ),
    .B1(\u_ppwm/u_mem/_0418_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0972_  (.B1(net434),
    .Y(\u_ppwm/u_mem/_0419_ ),
    .A1(net355),
    .A2(\u_ppwm/u_mem/memory[56] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0973_  (.A1(net355),
    .A2(\u_ppwm/u_mem/_0181_ ),
    .Y(\u_ppwm/u_mem/_0063_ ),
    .B1(\u_ppwm/u_mem/_0419_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0974_  (.B1(net434),
    .Y(\u_ppwm/u_mem/_0420_ ),
    .A1(net355),
    .A2(net214));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0975_  (.A1(net350),
    .A2(\u_ppwm/u_mem/_0180_ ),
    .Y(\u_ppwm/u_mem/_0064_ ),
    .B1(\u_ppwm/u_mem/_0420_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0976_  (.B1(net431),
    .Y(\u_ppwm/u_mem/_0421_ ),
    .A1(net351),
    .A2(net224));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0977_  (.A1(net349),
    .A2(\u_ppwm/u_mem/_0179_ ),
    .Y(\u_ppwm/u_mem/_0065_ ),
    .B1(\u_ppwm/u_mem/_0421_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0978_  (.B1(net430),
    .Y(\u_ppwm/u_mem/_0422_ ),
    .A1(net349),
    .A2(net253));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0979_  (.A1(net349),
    .A2(\u_ppwm/u_mem/_0178_ ),
    .Y(\u_ppwm/u_mem/_0066_ ),
    .B1(\u_ppwm/u_mem/_0422_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0980_  (.B1(net430),
    .Y(\u_ppwm/u_mem/_0423_ ),
    .A1(net348),
    .A2(\u_ppwm/u_mem/memory[60] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0981_  (.A1(net348),
    .A2(\u_ppwm/u_mem/_0177_ ),
    .Y(\u_ppwm/u_mem/_0067_ ),
    .B1(\u_ppwm/u_mem/_0423_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0982_  (.B1(net430),
    .Y(\u_ppwm/u_mem/_0424_ ),
    .A1(net348),
    .A2(net287));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0983_  (.A1(net348),
    .A2(\u_ppwm/u_mem/_0176_ ),
    .Y(\u_ppwm/u_mem/_0068_ ),
    .B1(\u_ppwm/u_mem/_0424_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0984_  (.B1(net431),
    .Y(\u_ppwm/u_mem/_0425_ ),
    .A1(net350),
    .A2(\u_ppwm/u_mem/memory[62] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0985_  (.A1(net351),
    .A2(\u_ppwm/u_mem/_0175_ ),
    .Y(\u_ppwm/u_mem/_0069_ ),
    .B1(\u_ppwm/u_mem/_0425_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0986_  (.B1(net434),
    .Y(\u_ppwm/u_mem/_0426_ ),
    .A1(net351),
    .A2(\u_ppwm/u_mem/memory[63] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0987_  (.A1(net351),
    .A2(\u_ppwm/u_mem/_0174_ ),
    .Y(\u_ppwm/u_mem/_0070_ ),
    .B1(\u_ppwm/u_mem/_0426_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0988_  (.B1(net431),
    .Y(\u_ppwm/u_mem/_0427_ ),
    .A1(net351),
    .A2(\u_ppwm/u_mem/memory[64] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0989_  (.A1(net351),
    .A2(\u_ppwm/u_mem/_0173_ ),
    .Y(\u_ppwm/u_mem/_0071_ ),
    .B1(\u_ppwm/u_mem/_0427_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0990_  (.B1(net431),
    .Y(\u_ppwm/u_mem/_0428_ ),
    .A1(net351),
    .A2(net270));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0991_  (.A1(net349),
    .A2(\u_ppwm/u_mem/_0172_ ),
    .Y(\u_ppwm/u_mem/_0072_ ),
    .B1(\u_ppwm/u_mem/_0428_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0992_  (.B1(net430),
    .Y(\u_ppwm/u_mem/_0429_ ),
    .A1(net349),
    .A2(\u_ppwm/u_mem/memory[66] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0993_  (.A1(net349),
    .A2(\u_ppwm/u_mem/_0171_ ),
    .Y(\u_ppwm/u_mem/_0073_ ),
    .B1(\u_ppwm/u_mem/_0429_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0994_  (.B1(net431),
    .Y(\u_ppwm/u_mem/_0430_ ),
    .A1(net348),
    .A2(\u_ppwm/u_mem/memory[67] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0995_  (.A1(net348),
    .A2(\u_ppwm/u_mem/_0170_ ),
    .Y(\u_ppwm/u_mem/_0074_ ),
    .B1(\u_ppwm/u_mem/_0430_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0996_  (.B1(net430),
    .Y(\u_ppwm/u_mem/_0431_ ),
    .A1(net346),
    .A2(net208));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0997_  (.A1(net346),
    .A2(\u_ppwm/u_mem/_0169_ ),
    .Y(\u_ppwm/u_mem/_0075_ ),
    .B1(\u_ppwm/u_mem/_0431_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_0998_  (.B1(net432),
    .Y(\u_ppwm/u_mem/_0432_ ),
    .A1(net350),
    .A2(\u_ppwm/u_mem/memory[69] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_0999_  (.A1(net350),
    .A2(\u_ppwm/u_mem/_0168_ ),
    .Y(\u_ppwm/u_mem/_0076_ ),
    .B1(\u_ppwm/u_mem/_0432_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1000_  (.B1(net434),
    .Y(\u_ppwm/u_mem/_0433_ ),
    .A1(net350),
    .A2(\u_ppwm/u_mem/memory[70] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1001_  (.A1(net350),
    .A2(\u_ppwm/u_mem/_0167_ ),
    .Y(\u_ppwm/u_mem/_0077_ ),
    .B1(\u_ppwm/u_mem/_0433_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1002_  (.B1(net434),
    .Y(\u_ppwm/u_mem/_0434_ ),
    .A1(net356),
    .A2(net276));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1003_  (.A1(net356),
    .A2(\u_ppwm/u_mem/_0166_ ),
    .Y(\u_ppwm/u_mem/_0078_ ),
    .B1(\u_ppwm/u_mem/_0434_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1004_  (.B1(net431),
    .Y(\u_ppwm/u_mem/_0435_ ),
    .A1(net350),
    .A2(net278));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1005_  (.A1(net350),
    .A2(\u_ppwm/u_mem/_0165_ ),
    .Y(\u_ppwm/u_mem/_0079_ ),
    .B1(\u_ppwm/u_mem/_0435_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1006_  (.B1(net431),
    .Y(\u_ppwm/u_mem/_0436_ ),
    .A1(net348),
    .A2(\u_ppwm/u_mem/memory[73] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1007_  (.A1(net348),
    .A2(\u_ppwm/u_mem/_0164_ ),
    .Y(\u_ppwm/u_mem/_0080_ ),
    .B1(\u_ppwm/u_mem/_0436_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1008_  (.B1(net430),
    .Y(\u_ppwm/u_mem/_0437_ ),
    .A1(net346),
    .A2(net293));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1009_  (.A1(net347),
    .A2(\u_ppwm/u_mem/_0163_ ),
    .Y(\u_ppwm/u_mem/_0081_ ),
    .B1(\u_ppwm/u_mem/_0437_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1010_  (.B1(net430),
    .Y(\u_ppwm/u_mem/_0438_ ),
    .A1(net346),
    .A2(net524));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1011_  (.A1(net346),
    .A2(\u_ppwm/u_mem/_0162_ ),
    .Y(\u_ppwm/u_mem/_0082_ ),
    .B1(\u_ppwm/u_mem/_0438_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1012_  (.B1(net429),
    .Y(\u_ppwm/u_mem/_0439_ ),
    .A1(net346),
    .A2(\u_ppwm/u_mem/memory[76] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1013_  (.A1(net357),
    .A2(\u_ppwm/u_mem/_0161_ ),
    .Y(\u_ppwm/u_mem/_0083_ ),
    .B1(\u_ppwm/u_mem/_0439_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1014_  (.B1(net434),
    .Y(\u_ppwm/u_mem/_0440_ ),
    .A1(net353),
    .A2(\u_ppwm/u_mem/memory[77] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1015_  (.A1(net355),
    .A2(\u_ppwm/u_mem/_0160_ ),
    .Y(\u_ppwm/u_mem/_0084_ ),
    .B1(\u_ppwm/u_mem/_0440_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1016_  (.B1(net435),
    .Y(\u_ppwm/u_mem/_0441_ ),
    .A1(net355),
    .A2(net229));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1017_  (.A1(net355),
    .A2(\u_ppwm/u_mem/_0159_ ),
    .Y(\u_ppwm/u_mem/_0085_ ),
    .B1(\u_ppwm/u_mem/_0441_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1018_  (.B1(net434),
    .Y(\u_ppwm/u_mem/_0442_ ),
    .A1(net355),
    .A2(\u_ppwm/u_mem/memory[79] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1019_  (.A1(net355),
    .A2(\u_ppwm/u_mem/_0158_ ),
    .Y(\u_ppwm/u_mem/_0086_ ),
    .B1(\u_ppwm/u_mem/_0442_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1020_  (.B1(net432),
    .Y(\u_ppwm/u_mem/_0443_ ),
    .A1(net347),
    .A2(\u_ppwm/u_mem/memory[80] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1021_  (.A1(net347),
    .A2(\u_ppwm/u_mem/_0157_ ),
    .Y(\u_ppwm/u_mem/_0087_ ),
    .B1(\u_ppwm/u_mem/_0443_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1022_  (.B1(net430),
    .Y(\u_ppwm/u_mem/_0444_ ),
    .A1(net347),
    .A2(\u_ppwm/u_mem/memory[81] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1023_  (.A1(net347),
    .A2(\u_ppwm/u_mem/_0156_ ),
    .Y(\u_ppwm/u_mem/_0088_ ),
    .B1(\u_ppwm/u_mem/_0444_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1024_  (.B1(net428),
    .Y(\u_ppwm/u_mem/_0445_ ),
    .A1(net346),
    .A2(net225));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1025_  (.A1(net346),
    .A2(\u_ppwm/u_mem/_0155_ ),
    .Y(\u_ppwm/u_mem/_0089_ ),
    .B1(\u_ppwm/u_mem/_0445_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1026_  (.B1(net428),
    .Y(\u_ppwm/u_mem/_0446_ ),
    .A1(net340),
    .A2(net516));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1027_  (.A1(net341),
    .A2(\u_ppwm/u_mem/_0154_ ),
    .Y(\u_ppwm/u_mem/_0090_ ),
    .B1(\u_ppwm/u_mem/_0446_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1028_  (.B1(net429),
    .Y(\u_ppwm/u_mem/_0447_ ),
    .A1(net347),
    .A2(\u_ppwm/u_mem/memory[84] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1029_  (.A1(net347),
    .A2(\u_ppwm/u_mem/_0153_ ),
    .Y(\u_ppwm/u_mem/_0091_ ),
    .B1(\u_ppwm/u_mem/_0447_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1030_  (.B1(net434),
    .Y(\u_ppwm/u_mem/_0448_ ),
    .A1(net353),
    .A2(\u_ppwm/u_mem/memory[85] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1031_  (.A1(net353),
    .A2(\u_ppwm/u_mem/_0152_ ),
    .Y(\u_ppwm/u_mem/_0092_ ),
    .B1(\u_ppwm/u_mem/_0448_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1032_  (.B1(net435),
    .Y(\u_ppwm/u_mem/_0449_ ),
    .A1(net353),
    .A2(net231));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1033_  (.A1(net353),
    .A2(\u_ppwm/u_mem/_0151_ ),
    .Y(\u_ppwm/u_mem/_0093_ ),
    .B1(\u_ppwm/u_mem/_0449_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1034_  (.B1(net433),
    .Y(\u_ppwm/u_mem/_0450_ ),
    .A1(net354),
    .A2(\u_ppwm/u_mem/memory[87] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1035_  (.A1(net354),
    .A2(\u_ppwm/u_mem/_0150_ ),
    .Y(\u_ppwm/u_mem/_0094_ ),
    .B1(\u_ppwm/u_mem/_0450_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1036_  (.B1(net433),
    .Y(\u_ppwm/u_mem/_0451_ ),
    .A1(net344),
    .A2(\u_ppwm/u_mem/memory[88] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1037_  (.A1(net344),
    .A2(\u_ppwm/u_mem/_0149_ ),
    .Y(\u_ppwm/u_mem/_0095_ ),
    .B1(\u_ppwm/u_mem/_0451_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1038_  (.B1(net433),
    .Y(\u_ppwm/u_mem/_0452_ ),
    .A1(net344),
    .A2(\u_ppwm/u_mem/memory[89] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1039_  (.A1(net344),
    .A2(\u_ppwm/u_mem/_0148_ ),
    .Y(\u_ppwm/u_mem/_0096_ ),
    .B1(\u_ppwm/u_mem/_0452_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1040_  (.B1(net433),
    .Y(\u_ppwm/u_mem/_0453_ ),
    .A1(net344),
    .A2(net210));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1041_  (.A1(net344),
    .A2(\u_ppwm/u_mem/_0147_ ),
    .Y(\u_ppwm/u_mem/_0097_ ),
    .B1(\u_ppwm/u_mem/_0453_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1042_  (.B1(net433),
    .Y(\u_ppwm/u_mem/_0454_ ),
    .A1(net342),
    .A2(net266));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1043_  (.A1(net342),
    .A2(\u_ppwm/u_mem/_0146_ ),
    .Y(\u_ppwm/u_mem/_0098_ ),
    .B1(\u_ppwm/u_mem/_0454_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1044_  (.B1(net433),
    .Y(\u_ppwm/u_mem/_0455_ ),
    .A1(net353),
    .A2(\u_ppwm/u_mem/memory[92] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1045_  (.A1(net353),
    .A2(\u_ppwm/u_mem/_0145_ ),
    .Y(\u_ppwm/u_mem/_0099_ ),
    .B1(\u_ppwm/u_mem/_0455_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1046_  (.B1(net435),
    .Y(\u_ppwm/u_mem/_0456_ ),
    .A1(net353),
    .A2(net274));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1047_  (.A1(net354),
    .A2(\u_ppwm/u_mem/_0144_ ),
    .Y(\u_ppwm/u_mem/_0100_ ),
    .B1(\u_ppwm/u_mem/_0456_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1048_  (.B1(net433),
    .Y(\u_ppwm/u_mem/_0457_ ),
    .A1(net354),
    .A2(\u_ppwm/u_mem/memory[94] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1049_  (.A1(net354),
    .A2(\u_ppwm/u_mem/_0143_ ),
    .Y(\u_ppwm/u_mem/_0101_ ),
    .B1(\u_ppwm/u_mem/_0457_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1050_  (.B1(net436),
    .Y(\u_ppwm/u_mem/_0458_ ),
    .A1(net345),
    .A2(net295));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1051_  (.A1(net345),
    .A2(\u_ppwm/u_mem/_0142_ ),
    .Y(\u_ppwm/u_mem/_0102_ ),
    .B1(\u_ppwm/u_mem/_0458_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1052_  (.B1(net433),
    .Y(\u_ppwm/u_mem/_0459_ ),
    .A1(net344),
    .A2(net473));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1053_  (.A1(net344),
    .A2(\u_ppwm/u_mem/_0141_ ),
    .Y(\u_ppwm/u_mem/_0103_ ),
    .B1(\u_ppwm/u_mem/_0459_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1054_  (.B1(net429),
    .Y(\u_ppwm/u_mem/_0460_ ),
    .A1(net342),
    .A2(\u_ppwm/u_mem/memory[97] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1055_  (.A1(net342),
    .A2(\u_ppwm/u_mem/_0140_ ),
    .Y(\u_ppwm/u_mem/_0104_ ),
    .B1(\u_ppwm/u_mem/_0460_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1056_  (.B1(net428),
    .Y(\u_ppwm/u_mem/_0461_ ),
    .A1(net341),
    .A2(\u_ppwm/u_mem/memory[98] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1057_  (.A1(net341),
    .A2(\u_ppwm/u_mem/_0139_ ),
    .Y(\u_ppwm/u_mem/_0105_ ),
    .B1(\u_ppwm/u_mem/_0461_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1058_  (.B1(net428),
    .Y(\u_ppwm/u_mem/_0462_ ),
    .A1(net341),
    .A2(net212));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1059_  (.A1(net341),
    .A2(\u_ppwm/u_mem/_0138_ ),
    .Y(\u_ppwm/u_mem/_0106_ ),
    .B1(\u_ppwm/u_mem/_0462_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1060_  (.B1(net428),
    .Y(\u_ppwm/u_mem/_0463_ ),
    .A1(net340),
    .A2(net286));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1061_  (.A1(net340),
    .A2(\u_ppwm/u_mem/_0137_ ),
    .Y(\u_ppwm/u_mem/_0107_ ),
    .B1(\u_ppwm/u_mem/_0463_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1062_  (.B1(net429),
    .Y(\u_ppwm/u_mem/_0464_ ),
    .A1(net342),
    .A2(\u_ppwm/u_mem/memory[101] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1063_  (.A1(net343),
    .A2(\u_ppwm/u_mem/_0136_ ),
    .Y(\u_ppwm/u_mem/_0108_ ),
    .B1(\u_ppwm/u_mem/_0464_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1064_  (.B1(net429),
    .Y(\u_ppwm/u_mem/_0465_ ),
    .A1(net339),
    .A2(net471));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1065_  (.A1(net339),
    .A2(\u_ppwm/u_mem/_0135_ ),
    .Y(\u_ppwm/u_mem/_0109_ ),
    .B1(\u_ppwm/u_mem/_0465_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1066_  (.B1(net423),
    .Y(\u_ppwm/u_mem/_0466_ ),
    .A1(net339),
    .A2(\u_ppwm/u_mem/memory[103] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1067_  (.A1(net339),
    .A2(\u_ppwm/u_mem/_0134_ ),
    .Y(\u_ppwm/u_mem/_0110_ ),
    .B1(\u_ppwm/u_mem/_0466_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1068_  (.B1(net429),
    .Y(\u_ppwm/u_mem/_0467_ ),
    .A1(net338),
    .A2(net477));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1069_  (.A1(net338),
    .A2(\u_ppwm/u_mem/_0133_ ),
    .Y(\u_ppwm/u_mem/_0111_ ),
    .B1(\u_ppwm/u_mem/_0467_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1070_  (.B1(net428),
    .Y(\u_ppwm/u_mem/_0468_ ),
    .A1(net340),
    .A2(\u_ppwm/u_mem/memory[105] ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1071_  (.A1(net338),
    .A2(\u_ppwm/u_mem/_0132_ ),
    .Y(\u_ppwm/u_mem/_0112_ ),
    .B1(\u_ppwm/u_mem/_0468_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1072_  (.B1(net428),
    .Y(\u_ppwm/u_mem/_0469_ ),
    .A1(net340),
    .A2(net233));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1073_  (.A1(net340),
    .A2(\u_ppwm/u_mem/_0131_ ),
    .Y(\u_ppwm/u_mem/_0113_ ),
    .B1(\u_ppwm/u_mem/_0469_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1074_  (.B1(net428),
    .Y(\u_ppwm/u_mem/_0470_ ),
    .A1(net340),
    .A2(net543));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1075_  (.A1(net340),
    .A2(\u_ppwm/u_mem/_0130_ ),
    .Y(\u_ppwm/u_mem/_0114_ ),
    .B1(\u_ppwm/u_mem/_0470_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1076_  (.B1(net429),
    .Y(\u_ppwm/u_mem/_0471_ ),
    .A1(net343),
    .A2(net558));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1077_  (.A1(net342),
    .A2(\u_ppwm/u_mem/_0129_ ),
    .Y(\u_ppwm/u_mem/_0115_ ),
    .B1(\u_ppwm/u_mem/_0471_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1078_  (.B1(net426),
    .Y(\u_ppwm/u_mem/_0472_ ),
    .A1(net345),
    .A2(\u_ppwm/u_mem/_0001_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1079_  (.A1(net345),
    .A2(\u_ppwm/u_mem/_0128_ ),
    .Y(\u_ppwm/u_mem/_0116_ ),
    .B1(\u_ppwm/u_mem/_0472_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1080_  (.B1(net426),
    .Y(\u_ppwm/u_mem/_0473_ ),
    .A1(net345),
    .A2(\u_ppwm/u_mem/_0002_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1081_  (.A1(\u_ppwm/u_mem/_0126_ ),
    .A2(net339),
    .Y(\u_ppwm/u_mem/_0117_ ),
    .B1(\u_ppwm/u_mem/_0473_ ));
 sg13g2_o21ai_1 \u_ppwm/u_mem/_1082_  (.B1(net423),
    .Y(\u_ppwm/u_mem/_0474_ ),
    .A1(net206),
    .A2(net339));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1083_  (.A1(\u_ppwm/u_mem/_0127_ ),
    .A2(net339),
    .Y(\u_ppwm/u_mem/_0118_ ),
    .B1(\u_ppwm/u_mem/_0474_ ));
 sg13g2_nand2b_2 \u_ppwm/u_mem/_1084_  (.Y(\u_ppwm/u_mem/_0475_ ),
    .B(net513),
    .A_N(net338));
 sg13g2_nand2_2 \u_ppwm/u_mem/_1085_  (.Y(\u_ppwm/u_mem/_0476_ ),
    .A(net423),
    .B(\u_ppwm/u_mem/_0475_ ));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1086_  (.A(net618),
    .B(net338),
    .Y(\u_ppwm/u_mem/_0477_ ));
 sg13g2_and2_1 \u_ppwm/u_mem/_1087_  (.A(net618),
    .B(net338),
    .X(\u_ppwm/u_mem/_0478_ ));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1088_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(\u_ppwm/u_mem/_0477_ ),
    .C(\u_ppwm/u_mem/_0478_ ),
    .Y(\u_ppwm/u_mem/_0119_ ));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1089_  (.A(net619),
    .B(\u_ppwm/u_mem/_0478_ ),
    .Y(\u_ppwm/u_mem/_0479_ ));
 sg13g2_and2_1 \u_ppwm/u_mem/_1090_  (.A(net619),
    .B(\u_ppwm/u_mem/_0478_ ),
    .X(\u_ppwm/u_mem/_0480_ ));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1091_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(\u_ppwm/u_mem/_0479_ ),
    .C(\u_ppwm/u_mem/_0480_ ),
    .Y(\u_ppwm/u_mem/_0120_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1092_  (.A1(net582),
    .A2(\u_ppwm/u_mem/_0475_ ),
    .Y(\u_ppwm/u_mem/_0481_ ),
    .B1(\u_ppwm/u_mem/_0480_ ));
 sg13g2_and4_1 \u_ppwm/u_mem/_1093_  (.A(net582),
    .B(net619),
    .C(net618),
    .D(net338),
    .X(\u_ppwm/u_mem/_0482_ ));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1094_  (.A(\u_ppwm/u_mem/_0238_ ),
    .B(net583),
    .C(\u_ppwm/u_mem/_0482_ ),
    .Y(\u_ppwm/u_mem/_0121_ ));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1095_  (.A(net624),
    .B(\u_ppwm/u_mem/_0482_ ),
    .Y(\u_ppwm/u_mem/_0483_ ));
 sg13g2_and2_1 \u_ppwm/u_mem/_1096_  (.A(net624),
    .B(\u_ppwm/u_mem/_0482_ ),
    .X(\u_ppwm/u_mem/_0484_ ));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1097_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(\u_ppwm/u_mem/_0483_ ),
    .C(\u_ppwm/u_mem/_0484_ ),
    .Y(\u_ppwm/u_mem/_0122_ ));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1098_  (.A(net602),
    .B(\u_ppwm/u_mem/_0484_ ),
    .Y(\u_ppwm/u_mem/_0485_ ));
 sg13g2_and3_1 \u_ppwm/u_mem/_1099_  (.X(\u_ppwm/u_mem/_0486_ ),
    .A(net602),
    .B(net624),
    .C(\u_ppwm/u_mem/_0482_ ));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1100_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(\u_ppwm/u_mem/_0485_ ),
    .C(\u_ppwm/u_mem/_0486_ ),
    .Y(\u_ppwm/u_mem/_0123_ ));
 sg13g2_nor2_1 \u_ppwm/u_mem/_1101_  (.A(net597),
    .B(\u_ppwm/u_mem/_0486_ ),
    .Y(\u_ppwm/u_mem/_0487_ ));
 sg13g2_and4_1 \u_ppwm/u_mem/_1102_  (.A(net597),
    .B(\u_ppwm/u_mem/bit_count[4] ),
    .C(\u_ppwm/u_mem/bit_count[3] ),
    .D(\u_ppwm/u_mem/_0482_ ),
    .X(\u_ppwm/u_mem/_0488_ ));
 sg13g2_nor3_1 \u_ppwm/u_mem/_1103_  (.A(\u_ppwm/u_mem/_0476_ ),
    .B(net598),
    .C(\u_ppwm/u_mem/_0488_ ),
    .Y(\u_ppwm/u_mem/_0124_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1104_  (.A1(net549),
    .A2(\u_ppwm/u_mem/_0475_ ),
    .Y(\u_ppwm/u_mem/_0489_ ),
    .B1(\u_ppwm/u_mem/_0488_ ));
 sg13g2_a21oi_1 \u_ppwm/u_mem/_1105_  (.A1(net549),
    .A2(\u_ppwm/u_mem/_0488_ ),
    .Y(\u_ppwm/u_mem/_0490_ ),
    .B1(\u_ppwm/u_mem/_0238_ ));
 sg13g2_nor2b_1 \u_ppwm/u_mem/_1106_  (.A(net550),
    .B_N(\u_ppwm/u_mem/_0490_ ),
    .Y(\u_ppwm/u_mem/_0125_ ));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1107_  (.RESET_B(net173),
    .D(net512),
    .Q(\u_ppwm/u_mem/memory[0] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1108_  (.RESET_B(net145),
    .D(\u_ppwm/u_mem/_0008_ ),
    .Q(\u_ppwm/u_mem/memory[1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1109_  (.RESET_B(net143),
    .D(net502),
    .Q(\u_ppwm/u_mem/memory[2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1110_  (.RESET_B(net141),
    .D(\u_ppwm/u_mem/_0010_ ),
    .Q(\u_ppwm/u_mem/memory[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1111_  (.RESET_B(net139),
    .D(net533),
    .Q(\u_ppwm/u_mem/memory[4] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1112_  (.RESET_B(net137),
    .D(net601),
    .Q(\u_ppwm/u_mem/memory[5] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1113_  (.RESET_B(net135),
    .D(net482),
    .Q(\u_ppwm/u_mem/memory[6] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1114_  (.RESET_B(net133),
    .D(net561),
    .Q(\u_ppwm/u_mem/memory[7] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1115_  (.RESET_B(net131),
    .D(net242),
    .Q(\u_ppwm/u_mem/memory[8] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1116_  (.RESET_B(net129),
    .D(\u_ppwm/u_mem/_0016_ ),
    .Q(\u_ppwm/u_mem/memory[9] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1117_  (.RESET_B(net127),
    .D(net465),
    .Q(\u_ppwm/u_mem/memory[10] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1118_  (.RESET_B(net125),
    .D(net470),
    .Q(\u_ppwm/u_mem/memory[11] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1119_  (.RESET_B(net123),
    .D(net492),
    .Q(\u_ppwm/u_mem/memory[12] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1120_  (.RESET_B(net121),
    .D(net507),
    .Q(\u_ppwm/u_mem/memory[13] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1121_  (.RESET_B(net119),
    .D(net590),
    .Q(\u_ppwm/u_mem/memory[14] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1122_  (.RESET_B(net117),
    .D(\u_ppwm/u_mem/_0022_ ),
    .Q(\u_ppwm/u_mem/memory[15] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1123_  (.RESET_B(net115),
    .D(net484),
    .Q(\u_ppwm/u_mem/memory[16] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1124_  (.RESET_B(net113),
    .D(net302),
    .Q(\u_ppwm/u_mem/memory[17] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1125_  (.RESET_B(net111),
    .D(net504),
    .Q(\u_ppwm/u_mem/memory[18] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1126_  (.RESET_B(net109),
    .D(\u_ppwm/u_mem/_0026_ ),
    .Q(\u_ppwm/u_mem/memory[19] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1127_  (.RESET_B(net107),
    .D(net480),
    .Q(\u_ppwm/u_mem/memory[20] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1128_  (.RESET_B(net105),
    .D(\u_ppwm/u_mem/_0028_ ),
    .Q(\u_ppwm/u_mem/memory[21] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1129_  (.RESET_B(net103),
    .D(\u_ppwm/u_mem/_0029_ ),
    .Q(\u_ppwm/u_mem/memory[22] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1130_  (.RESET_B(net101),
    .D(net476),
    .Q(\u_ppwm/u_mem/memory[23] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1131_  (.RESET_B(net99),
    .D(net300),
    .Q(\u_ppwm/u_mem/memory[24] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1132_  (.RESET_B(net97),
    .D(net571),
    .Q(\u_ppwm/u_mem/memory[25] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1133_  (.RESET_B(net95),
    .D(net255),
    .Q(\u_ppwm/u_mem/memory[26] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1134_  (.RESET_B(net93),
    .D(net236),
    .Q(\u_ppwm/u_mem/memory[27] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1135_  (.RESET_B(net91),
    .D(\u_ppwm/u_mem/_0035_ ),
    .Q(\u_ppwm/u_mem/memory[28] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1136_  (.RESET_B(net89),
    .D(net531),
    .Q(\u_ppwm/u_mem/memory[29] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1137_  (.RESET_B(net87),
    .D(net518),
    .Q(\u_ppwm/u_mem/memory[30] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1138_  (.RESET_B(net85),
    .D(net217),
    .Q(\u_ppwm/u_mem/memory[31] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1139_  (.RESET_B(net83),
    .D(net273),
    .Q(\u_ppwm/u_mem/memory[32] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1140_  (.RESET_B(net81),
    .D(\u_ppwm/u_mem/_0040_ ),
    .Q(\u_ppwm/u_mem/memory[33] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1141_  (.RESET_B(net79),
    .D(net290),
    .Q(\u_ppwm/u_mem/memory[34] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1142_  (.RESET_B(net77),
    .D(net495),
    .Q(\u_ppwm/u_mem/memory[35] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1143_  (.RESET_B(net75),
    .D(net460),
    .Q(\u_ppwm/u_mem/memory[36] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1144_  (.RESET_B(net73),
    .D(\u_ppwm/u_mem/_0044_ ),
    .Q(\u_ppwm/u_mem/memory[37] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1145_  (.RESET_B(net71),
    .D(net281),
    .Q(\u_ppwm/u_mem/memory[38] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1146_  (.RESET_B(net69),
    .D(\u_ppwm/u_mem/_0046_ ),
    .Q(\u_ppwm/u_mem/memory[39] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1147_  (.RESET_B(net67),
    .D(net542),
    .Q(\u_ppwm/u_mem/memory[40] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1148_  (.RESET_B(net65),
    .D(net540),
    .Q(\u_ppwm/u_mem/memory[41] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1149_  (.RESET_B(net63),
    .D(net520),
    .Q(\u_ppwm/u_mem/memory[42] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1150_  (.RESET_B(net61),
    .D(\u_ppwm/u_mem/_0050_ ),
    .Q(\u_ppwm/u_mem/memory[43] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1151_  (.RESET_B(net59),
    .D(net298),
    .Q(\u_ppwm/u_mem/memory[44] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1152_  (.RESET_B(net57),
    .D(\u_ppwm/u_mem/_0052_ ),
    .Q(\u_ppwm/u_mem/memory[45] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1153_  (.RESET_B(net55),
    .D(net456),
    .Q(\u_ppwm/u_mem/memory[46] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1154_  (.RESET_B(net172),
    .D(net248),
    .Q(\u_ppwm/u_mem/memory[47] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1155_  (.RESET_B(net170),
    .D(\u_ppwm/u_mem/_0055_ ),
    .Q(\u_ppwm/u_mem/memory[48] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1156_  (.RESET_B(net168),
    .D(net261),
    .Q(\u_ppwm/u_mem/memory[49] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1157_  (.RESET_B(net166),
    .D(net238),
    .Q(\u_ppwm/u_mem/memory[50] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1158_  (.RESET_B(net164),
    .D(\u_ppwm/u_mem/_0058_ ),
    .Q(\u_ppwm/u_mem/memory[51] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1159_  (.RESET_B(net162),
    .D(\u_ppwm/u_mem/_0059_ ),
    .Q(\u_ppwm/u_mem/memory[52] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1160_  (.RESET_B(net160),
    .D(net257),
    .Q(\u_ppwm/u_mem/memory[53] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1161_  (.RESET_B(net158),
    .D(\u_ppwm/u_mem/_0061_ ),
    .Q(\u_ppwm/u_mem/memory[54] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1162_  (.RESET_B(net156),
    .D(net283),
    .Q(\u_ppwm/u_mem/memory[55] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1163_  (.RESET_B(net154),
    .D(net215),
    .Q(\u_ppwm/u_mem/memory[56] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1164_  (.RESET_B(net152),
    .D(\u_ppwm/u_mem/_0064_ ),
    .Q(\u_ppwm/u_mem/memory[57] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1165_  (.RESET_B(net150),
    .D(\u_ppwm/u_mem/_0065_ ),
    .Q(\u_ppwm/u_mem/memory[58] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1166_  (.RESET_B(net148),
    .D(\u_ppwm/u_mem/_0066_ ),
    .Q(\u_ppwm/u_mem/memory[59] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1167_  (.RESET_B(net146),
    .D(net288),
    .Q(\u_ppwm/u_mem/memory[60] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1168_  (.RESET_B(net142),
    .D(\u_ppwm/u_mem/_0068_ ),
    .Q(\u_ppwm/u_mem/memory[61] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1169_  (.RESET_B(net138),
    .D(net488),
    .Q(\u_ppwm/u_mem/memory[62] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1170_  (.RESET_B(net134),
    .D(net468),
    .Q(\u_ppwm/u_mem/memory[63] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1171_  (.RESET_B(net130),
    .D(net271),
    .Q(\u_ppwm/u_mem/memory[64] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1172_  (.RESET_B(net126),
    .D(\u_ppwm/u_mem/_0072_ ),
    .Q(\u_ppwm/u_mem/memory[65] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1173_  (.RESET_B(net122),
    .D(net244),
    .Q(\u_ppwm/u_mem/memory[66] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1174_  (.RESET_B(net118),
    .D(net209),
    .Q(\u_ppwm/u_mem/memory[67] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1175_  (.RESET_B(net114),
    .D(\u_ppwm/u_mem/_0075_ ),
    .Q(\u_ppwm/u_mem/memory[68] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1176_  (.RESET_B(net110),
    .D(net454),
    .Q(\u_ppwm/u_mem/memory[69] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1177_  (.RESET_B(net106),
    .D(net277),
    .Q(\u_ppwm/u_mem/memory[70] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1178_  (.RESET_B(net102),
    .D(net279),
    .Q(\u_ppwm/u_mem/memory[71] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1179_  (.RESET_B(net98),
    .D(\u_ppwm/u_mem/_0079_ ),
    .Q(\u_ppwm/u_mem/memory[72] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1180_  (.RESET_B(net94),
    .D(net294),
    .Q(\u_ppwm/u_mem/memory[73] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1181_  (.RESET_B(net90),
    .D(\u_ppwm/u_mem/_0081_ ),
    .Q(\u_ppwm/u_mem/memory[74] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1182_  (.RESET_B(net86),
    .D(\u_ppwm/u_mem/_0082_ ),
    .Q(\u_ppwm/u_mem/memory[75] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1183_  (.RESET_B(net82),
    .D(net526),
    .Q(\u_ppwm/u_mem/memory[76] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1184_  (.RESET_B(net78),
    .D(net230),
    .Q(\u_ppwm/u_mem/memory[77] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1185_  (.RESET_B(net74),
    .D(\u_ppwm/u_mem/_0085_ ),
    .Q(\u_ppwm/u_mem/memory[78] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1186_  (.RESET_B(net70),
    .D(net509),
    .Q(\u_ppwm/u_mem/memory[79] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1187_  (.RESET_B(net66),
    .D(net240),
    .Q(\u_ppwm/u_mem/memory[80] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1188_  (.RESET_B(net62),
    .D(net226),
    .Q(\u_ppwm/u_mem/memory[81] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1189_  (.RESET_B(net58),
    .D(\u_ppwm/u_mem/_0089_ ),
    .Q(\u_ppwm/u_mem/memory[82] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1190_  (.RESET_B(net54),
    .D(\u_ppwm/u_mem/_0090_ ),
    .Q(\u_ppwm/u_mem/memory[83] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1191_  (.RESET_B(net169),
    .D(net486),
    .Q(\u_ppwm/u_mem/memory[84] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1192_  (.RESET_B(net165),
    .D(net232),
    .Q(\u_ppwm/u_mem/memory[85] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1193_  (.RESET_B(net161),
    .D(net285),
    .Q(\u_ppwm/u_mem/memory[86] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1194_  (.RESET_B(net157),
    .D(net259),
    .Q(\u_ppwm/u_mem/memory[87] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1195_  (.RESET_B(net153),
    .D(net246),
    .Q(\u_ppwm/u_mem/memory[88] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1196_  (.RESET_B(net149),
    .D(net211),
    .Q(\u_ppwm/u_mem/memory[89] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1197_  (.RESET_B(net144),
    .D(net267),
    .Q(\u_ppwm/u_mem/memory[90] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1198_  (.RESET_B(net136),
    .D(net499),
    .Q(\u_ppwm/u_mem/memory[91] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1199_  (.RESET_B(net128),
    .D(net275),
    .Q(\u_ppwm/u_mem/memory[92] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1200_  (.RESET_B(net120),
    .D(\u_ppwm/u_mem/_0100_ ),
    .Q(\u_ppwm/u_mem/memory[93] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1201_  (.RESET_B(net112),
    .D(net296),
    .Q(\u_ppwm/u_mem/memory[94] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1202_  (.RESET_B(net104),
    .D(net474),
    .Q(\u_ppwm/u_mem/memory[95] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1203_  (.RESET_B(net96),
    .D(net490),
    .Q(\u_ppwm/u_mem/memory[96] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1204_  (.RESET_B(net88),
    .D(net263),
    .Q(\u_ppwm/u_mem/memory[97] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1205_  (.RESET_B(net80),
    .D(net213),
    .Q(\u_ppwm/u_mem/memory[98] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1206_  (.RESET_B(net72),
    .D(\u_ppwm/u_mem/_0106_ ),
    .Q(\u_ppwm/u_mem/memory[99] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1207_  (.RESET_B(net64),
    .D(\u_ppwm/u_mem/_0107_ ),
    .Q(\u_ppwm/u_mem/memory[100] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1208_  (.RESET_B(net56),
    .D(net472),
    .Q(\u_ppwm/u_mem/memory[101] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1209_  (.RESET_B(net167),
    .D(\u_ppwm/u_mem/_0109_ ),
    .Q(\u_ppwm/u_mem/memory[102] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1210_  (.RESET_B(net159),
    .D(net478),
    .Q(\u_ppwm/u_mem/memory[103] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1211_  (.RESET_B(net151),
    .D(net567),
    .Q(\u_ppwm/u_mem/memory[104] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1212_  (.RESET_B(net140),
    .D(net234),
    .Q(\u_ppwm/u_mem/memory[105] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1213_  (.RESET_B(net124),
    .D(\u_ppwm/u_mem/_0113_ ),
    .Q(\u_ppwm/u_mem/memory[106] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1214_  (.RESET_B(net108),
    .D(\u_ppwm/u_mem/_0114_ ),
    .Q(\u_ppwm/u_mem/memory[107] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1215_  (.RESET_B(net92),
    .D(net593),
    .Q(\u_ppwm/u_mem/_0000_ ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1216_  (.RESET_B(net76),
    .D(net522),
    .Q(\u_ppwm/u_mem/_0001_ ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1217_  (.RESET_B(net60),
    .D(net207),
    .Q(\u_ppwm/u_mem/_0002_ ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1218_  (.RESET_B(net163),
    .D(\u_ppwm/u_mem/_0118_ ),
    .Q(\u_ppwm/u_mem/_0003_ ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1219_  (.RESET_B(net147),
    .D(\u_ppwm/u_mem/_0119_ ),
    .Q(\u_ppwm/u_mem/bit_count[0] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1220_  (.RESET_B(net116),
    .D(\u_ppwm/u_mem/_0120_ ),
    .Q(\u_ppwm/u_mem/bit_count[1] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1221_  (.RESET_B(net84),
    .D(net584),
    .Q(\u_ppwm/u_mem/bit_count[2] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1222_  (.RESET_B(net171),
    .D(\u_ppwm/u_mem/_0122_ ),
    .Q(\u_ppwm/u_mem/bit_count[3] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1223_  (.RESET_B(net132),
    .D(\u_ppwm/u_mem/_0123_ ),
    .Q(\u_ppwm/u_mem/bit_count[4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1224_  (.RESET_B(net68),
    .D(net599),
    .Q(\u_ppwm/u_mem/bit_count[5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1225_  (.RESET_B(net174),
    .D(net551),
    .Q(\u_ppwm/u_mem/bit_count[6] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1226_  (.RESET_B(net175),
    .D(net514),
    .Q(\u_ppwm/u_mem/state_q[0] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_mem/_1227_  (.RESET_B(net155),
    .D(\u_ppwm/u_mem/_0005_ ),
    .Q(\u_ppwm/mem_write_done ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_mem/_1228_  (.RESET_B(net100),
    .D(\u_ppwm/u_mem/_0006_ ),
    .Q(\u_ppwm/u_mem/state_q[2] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_tiehi \u_ppwm/u_mem/_1153__55  (.L_HI(net55));
 sg13g2_tiehi \u_ppwm/u_mem/_1208__56  (.L_HI(net56));
 sg13g2_tiehi \u_ppwm/u_mem/_1152__57  (.L_HI(net57));
 sg13g2_tiehi \u_ppwm/u_mem/_1189__58  (.L_HI(net58));
 sg13g2_tiehi \u_ppwm/u_mem/_1151__59  (.L_HI(net59));
 sg13g2_tiehi \u_ppwm/u_mem/_1217__60  (.L_HI(net60));
 sg13g2_tiehi \u_ppwm/u_mem/_1150__61  (.L_HI(net61));
 sg13g2_tiehi \u_ppwm/u_mem/_1188__62  (.L_HI(net62));
 sg13g2_tiehi \u_ppwm/u_mem/_1149__63  (.L_HI(net63));
 sg13g2_tiehi \u_ppwm/u_mem/_1207__64  (.L_HI(net64));
 sg13g2_tiehi \u_ppwm/u_mem/_1148__65  (.L_HI(net65));
 sg13g2_tiehi \u_ppwm/u_mem/_1187__66  (.L_HI(net66));
 sg13g2_tiehi \u_ppwm/u_mem/_1147__67  (.L_HI(net67));
 sg13g2_tiehi \u_ppwm/u_mem/_1224__68  (.L_HI(net68));
 sg13g2_tiehi \u_ppwm/u_mem/_1146__69  (.L_HI(net69));
 sg13g2_tiehi \u_ppwm/u_mem/_1186__70  (.L_HI(net70));
 sg13g2_tiehi \u_ppwm/u_mem/_1145__71  (.L_HI(net71));
 sg13g2_tiehi \u_ppwm/u_mem/_1206__72  (.L_HI(net72));
 sg13g2_tiehi \u_ppwm/u_mem/_1144__73  (.L_HI(net73));
 sg13g2_tiehi \u_ppwm/u_mem/_1185__74  (.L_HI(net74));
 sg13g2_tiehi \u_ppwm/u_mem/_1143__75  (.L_HI(net75));
 sg13g2_tiehi \u_ppwm/u_mem/_1216__76  (.L_HI(net76));
 sg13g2_tiehi \u_ppwm/u_mem/_1142__77  (.L_HI(net77));
 sg13g2_tiehi \u_ppwm/u_mem/_1184__78  (.L_HI(net78));
 sg13g2_tiehi \u_ppwm/u_mem/_1141__79  (.L_HI(net79));
 sg13g2_tiehi \u_ppwm/u_mem/_1205__80  (.L_HI(net80));
 sg13g2_tiehi \u_ppwm/u_mem/_1140__81  (.L_HI(net81));
 sg13g2_tiehi \u_ppwm/u_mem/_1183__82  (.L_HI(net82));
 sg13g2_tiehi \u_ppwm/u_mem/_1139__83  (.L_HI(net83));
 sg13g2_tiehi \u_ppwm/u_mem/_1221__84  (.L_HI(net84));
 sg13g2_tiehi \u_ppwm/u_mem/_1138__85  (.L_HI(net85));
 sg13g2_tiehi \u_ppwm/u_mem/_1182__86  (.L_HI(net86));
 sg13g2_tiehi \u_ppwm/u_mem/_1137__87  (.L_HI(net87));
 sg13g2_tiehi \u_ppwm/u_mem/_1204__88  (.L_HI(net88));
 sg13g2_tiehi \u_ppwm/u_mem/_1136__89  (.L_HI(net89));
 sg13g2_tiehi \u_ppwm/u_mem/_1181__90  (.L_HI(net90));
 sg13g2_tiehi \u_ppwm/u_mem/_1135__91  (.L_HI(net91));
 sg13g2_tiehi \u_ppwm/u_mem/_1215__92  (.L_HI(net92));
 sg13g2_tiehi \u_ppwm/u_mem/_1134__93  (.L_HI(net93));
 sg13g2_tiehi \u_ppwm/u_mem/_1180__94  (.L_HI(net94));
 sg13g2_tiehi \u_ppwm/u_mem/_1133__95  (.L_HI(net95));
 sg13g2_tiehi \u_ppwm/u_mem/_1203__96  (.L_HI(net96));
 sg13g2_tiehi \u_ppwm/u_mem/_1132__97  (.L_HI(net97));
 sg13g2_tiehi \u_ppwm/u_mem/_1179__98  (.L_HI(net98));
 sg13g2_tiehi \u_ppwm/u_mem/_1131__99  (.L_HI(net99));
 sg13g2_tiehi \u_ppwm/u_mem/_1228__100  (.L_HI(net100));
 sg13g2_tiehi \u_ppwm/u_mem/_1130__101  (.L_HI(net101));
 sg13g2_tiehi \u_ppwm/u_mem/_1178__102  (.L_HI(net102));
 sg13g2_tiehi \u_ppwm/u_mem/_1129__103  (.L_HI(net103));
 sg13g2_tiehi \u_ppwm/u_mem/_1202__104  (.L_HI(net104));
 sg13g2_tiehi \u_ppwm/u_mem/_1128__105  (.L_HI(net105));
 sg13g2_tiehi \u_ppwm/u_mem/_1177__106  (.L_HI(net106));
 sg13g2_tiehi \u_ppwm/u_mem/_1127__107  (.L_HI(net107));
 sg13g2_tiehi \u_ppwm/u_mem/_1214__108  (.L_HI(net108));
 sg13g2_tiehi \u_ppwm/u_mem/_1126__109  (.L_HI(net109));
 sg13g2_tiehi \u_ppwm/u_mem/_1176__110  (.L_HI(net110));
 sg13g2_tiehi \u_ppwm/u_mem/_1125__111  (.L_HI(net111));
 sg13g2_tiehi \u_ppwm/u_mem/_1201__112  (.L_HI(net112));
 sg13g2_tiehi \u_ppwm/u_mem/_1124__113  (.L_HI(net113));
 sg13g2_tiehi \u_ppwm/u_mem/_1175__114  (.L_HI(net114));
 sg13g2_tiehi \u_ppwm/u_mem/_1123__115  (.L_HI(net115));
 sg13g2_tiehi \u_ppwm/u_mem/_1220__116  (.L_HI(net116));
 sg13g2_tiehi \u_ppwm/u_mem/_1122__117  (.L_HI(net117));
 sg13g2_tiehi \u_ppwm/u_mem/_1174__118  (.L_HI(net118));
 sg13g2_tiehi \u_ppwm/u_mem/_1121__119  (.L_HI(net119));
 sg13g2_tiehi \u_ppwm/u_mem/_1200__120  (.L_HI(net120));
 sg13g2_tiehi \u_ppwm/u_mem/_1120__121  (.L_HI(net121));
 sg13g2_tiehi \u_ppwm/u_mem/_1173__122  (.L_HI(net122));
 sg13g2_tiehi \u_ppwm/u_mem/_1119__123  (.L_HI(net123));
 sg13g2_tiehi \u_ppwm/u_mem/_1213__124  (.L_HI(net124));
 sg13g2_tiehi \u_ppwm/u_mem/_1118__125  (.L_HI(net125));
 sg13g2_tiehi \u_ppwm/u_mem/_1172__126  (.L_HI(net126));
 sg13g2_tiehi \u_ppwm/u_mem/_1117__127  (.L_HI(net127));
 sg13g2_tiehi \u_ppwm/u_mem/_1199__128  (.L_HI(net128));
 sg13g2_tiehi \u_ppwm/u_mem/_1116__129  (.L_HI(net129));
 sg13g2_tiehi \u_ppwm/u_mem/_1171__130  (.L_HI(net130));
 sg13g2_tiehi \u_ppwm/u_mem/_1115__131  (.L_HI(net131));
 sg13g2_tiehi \u_ppwm/u_mem/_1223__132  (.L_HI(net132));
 sg13g2_tiehi \u_ppwm/u_mem/_1114__133  (.L_HI(net133));
 sg13g2_tiehi \u_ppwm/u_mem/_1170__134  (.L_HI(net134));
 sg13g2_tiehi \u_ppwm/u_mem/_1113__135  (.L_HI(net135));
 sg13g2_tiehi \u_ppwm/u_mem/_1198__136  (.L_HI(net136));
 sg13g2_tiehi \u_ppwm/u_mem/_1112__137  (.L_HI(net137));
 sg13g2_tiehi \u_ppwm/u_mem/_1169__138  (.L_HI(net138));
 sg13g2_tiehi \u_ppwm/u_mem/_1111__139  (.L_HI(net139));
 sg13g2_tiehi \u_ppwm/u_mem/_1212__140  (.L_HI(net140));
 sg13g2_tiehi \u_ppwm/u_mem/_1110__141  (.L_HI(net141));
 sg13g2_tiehi \u_ppwm/u_mem/_1168__142  (.L_HI(net142));
 sg13g2_tiehi \u_ppwm/u_mem/_1109__143  (.L_HI(net143));
 sg13g2_tiehi \u_ppwm/u_mem/_1197__144  (.L_HI(net144));
 sg13g2_tiehi \u_ppwm/u_mem/_1108__145  (.L_HI(net145));
 sg13g2_tiehi \u_ppwm/u_mem/_1167__146  (.L_HI(net146));
 sg13g2_tiehi \u_ppwm/u_mem/_1219__147  (.L_HI(net147));
 sg13g2_tiehi \u_ppwm/u_mem/_1166__148  (.L_HI(net148));
 sg13g2_tiehi \u_ppwm/u_mem/_1196__149  (.L_HI(net149));
 sg13g2_tiehi \u_ppwm/u_mem/_1165__150  (.L_HI(net150));
 sg13g2_tiehi \u_ppwm/u_mem/_1211__151  (.L_HI(net151));
 sg13g2_tiehi \u_ppwm/u_mem/_1164__152  (.L_HI(net152));
 sg13g2_tiehi \u_ppwm/u_mem/_1195__153  (.L_HI(net153));
 sg13g2_tiehi \u_ppwm/u_mem/_1163__154  (.L_HI(net154));
 sg13g2_tiehi \u_ppwm/u_mem/_1227__155  (.L_HI(net155));
 sg13g2_tiehi \u_ppwm/u_mem/_1162__156  (.L_HI(net156));
 sg13g2_tiehi \u_ppwm/u_mem/_1194__157  (.L_HI(net157));
 sg13g2_tiehi \u_ppwm/u_mem/_1161__158  (.L_HI(net158));
 sg13g2_tiehi \u_ppwm/u_mem/_1210__159  (.L_HI(net159));
 sg13g2_tiehi \u_ppwm/u_mem/_1160__160  (.L_HI(net160));
 sg13g2_tiehi \u_ppwm/u_mem/_1193__161  (.L_HI(net161));
 sg13g2_tiehi \u_ppwm/u_mem/_1159__162  (.L_HI(net162));
 sg13g2_tiehi \u_ppwm/u_mem/_1218__163  (.L_HI(net163));
 sg13g2_tiehi \u_ppwm/u_mem/_1158__164  (.L_HI(net164));
 sg13g2_tiehi \u_ppwm/u_mem/_1192__165  (.L_HI(net165));
 sg13g2_tiehi \u_ppwm/u_mem/_1157__166  (.L_HI(net166));
 sg13g2_tiehi \u_ppwm/u_mem/_1209__167  (.L_HI(net167));
 sg13g2_tiehi \u_ppwm/u_mem/_1156__168  (.L_HI(net168));
 sg13g2_tiehi \u_ppwm/u_mem/_1191__169  (.L_HI(net169));
 sg13g2_tiehi \u_ppwm/u_mem/_1155__170  (.L_HI(net170));
 sg13g2_tiehi \u_ppwm/u_mem/_1222__171  (.L_HI(net171));
 sg13g2_tiehi \u_ppwm/u_mem/_1154__172  (.L_HI(net172));
 sg13g2_tiehi \u_ppwm/u_mem/_1107__173  (.L_HI(net173));
 sg13g2_tiehi \u_ppwm/u_mem/_1225__174  (.L_HI(net174));
 sg13g2_tiehi \u_ppwm/u_mem/_1226__175  (.L_HI(net175));
 sg13g2_tiehi \u_ppwm/u_pwm/_247__176  (.L_HI(net176));
 sg13g2_inv_2 \u_ppwm/u_pwm/_124_  (.Y(\u_ppwm/u_pwm/_069_ ),
    .A(net594));
 sg13g2_inv_2 \u_ppwm/u_pwm/_125_  (.Y(\u_ppwm/u_pwm/_070_ ),
    .A(net604));
 sg13g2_inv_1 \u_ppwm/u_pwm/_126_  (.Y(\u_ppwm/u_pwm/_071_ ),
    .A(net580));
 sg13g2_inv_1 \u_ppwm/u_pwm/_127_  (.Y(\u_ppwm/u_pwm/_072_ ),
    .A(\u_ppwm/u_pwm/counter[2] ));
 sg13g2_inv_1 \u_ppwm/u_pwm/_128_  (.Y(\u_ppwm/u_pwm/_073_ ),
    .A(\u_ppwm/u_pwm/counter[1] ));
 sg13g2_inv_1 \u_ppwm/u_pwm/_129_  (.Y(\u_ppwm/u_pwm/_074_ ),
    .A(net568));
 sg13g2_inv_1 \u_ppwm/u_pwm/_130_  (.Y(\u_ppwm/u_pwm/_075_ ),
    .A(net264));
 sg13g2_inv_1 \u_ppwm/u_pwm/_131_  (.Y(\u_ppwm/u_pwm/_076_ ),
    .A(net249));
 sg13g2_inv_1 \u_ppwm/u_pwm/_132_  (.Y(\u_ppwm/u_pwm/_077_ ),
    .A(net220));
 sg13g2_inv_1 \u_ppwm/u_pwm/_133_  (.Y(\u_ppwm/u_pwm/_078_ ),
    .A(net222));
 sg13g2_inv_1 \u_ppwm/u_pwm/_134_  (.Y(\u_ppwm/u_pwm/_079_ ),
    .A(net304));
 sg13g2_inv_1 \u_ppwm/u_pwm/_135_  (.Y(\u_ppwm/u_pwm/_080_ ),
    .A(net496));
 sg13g2_inv_1 \u_ppwm/u_pwm/_136_  (.Y(\u_ppwm/u_pwm/_081_ ),
    .A(net562));
 sg13g2_inv_1 \u_ppwm/u_pwm/_137_  (.Y(\u_ppwm/u_pwm/_082_ ),
    .A(net218));
 sg13g2_inv_1 \u_ppwm/u_pwm/_138_  (.Y(\u_ppwm/u_pwm/_083_ ),
    .A(net200));
 sg13g2_inv_1 \u_ppwm/u_pwm/_139_  (.Y(\u_ppwm/u_pwm/_084_ ),
    .A(net422));
 sg13g2_nor4_1 \u_ppwm/u_pwm/_140_  (.A(net337),
    .B(\u_ppwm/u_pwm/counter[2] ),
    .C(\u_ppwm/u_pwm/counter[1] ),
    .D(\u_ppwm/u_pwm/counter[0] ),
    .Y(\u_ppwm/u_pwm/_085_ ));
 sg13g2_nor4_1 \u_ppwm/u_pwm/_141_  (.A(\u_ppwm/u_pwm/counter[7] ),
    .B(\u_ppwm/u_pwm/counter[6] ),
    .C(\u_ppwm/u_pwm/counter[5] ),
    .D(\u_ppwm/u_pwm/counter[4] ),
    .Y(\u_ppwm/u_pwm/_086_ ));
 sg13g2_nand4_1 \u_ppwm/u_pwm/_142_  (.B(\u_ppwm/u_pwm/_070_ ),
    .C(\u_ppwm/u_pwm/_085_ ),
    .A(\u_ppwm/u_pwm/_069_ ),
    .Y(\u_ppwm/u_pwm/_087_ ),
    .D(\u_ppwm/u_pwm/_086_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_143_  (.B1(net424),
    .Y(\u_ppwm/u_pwm/_088_ ),
    .A1(\u_ppwm/pwm_value[0] ),
    .A2(net328));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_144_  (.A1(\u_ppwm/u_pwm/_083_ ),
    .A2(net328),
    .Y(\u_ppwm/u_pwm/_000_ ),
    .B1(\u_ppwm/u_pwm/_088_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_145_  (.B1(net424),
    .Y(\u_ppwm/u_pwm/_089_ ),
    .A1(net398),
    .A2(net328));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_146_  (.A1(\u_ppwm/u_pwm/_082_ ),
    .A2(net328),
    .Y(\u_ppwm/u_pwm/_001_ ),
    .B1(\u_ppwm/u_pwm/_089_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_147_  (.B1(net425),
    .Y(\u_ppwm/u_pwm/_090_ ),
    .A1(net396),
    .A2(net329));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_148_  (.A1(\u_ppwm/u_pwm/_081_ ),
    .A2(net328),
    .Y(\u_ppwm/u_pwm/_002_ ),
    .B1(\u_ppwm/u_pwm/_090_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_149_  (.B1(net424),
    .Y(\u_ppwm/u_pwm/_091_ ),
    .A1(net394),
    .A2(net329));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_150_  (.A1(\u_ppwm/u_pwm/_080_ ),
    .A2(net328),
    .Y(\u_ppwm/u_pwm/_003_ ),
    .B1(\u_ppwm/u_pwm/_091_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_151_  (.B1(net425),
    .Y(\u_ppwm/u_pwm/_092_ ),
    .A1(net392),
    .A2(net330));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_152_  (.A1(\u_ppwm/u_pwm/_079_ ),
    .A2(net330),
    .Y(\u_ppwm/u_pwm/_004_ ),
    .B1(\u_ppwm/u_pwm/_092_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_153_  (.B1(net424),
    .Y(\u_ppwm/u_pwm/_093_ ),
    .A1(net391),
    .A2(net330));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_154_  (.A1(\u_ppwm/u_pwm/_078_ ),
    .A2(net330),
    .Y(\u_ppwm/u_pwm/_005_ ),
    .B1(\u_ppwm/u_pwm/_093_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_155_  (.B1(net424),
    .Y(\u_ppwm/u_pwm/_094_ ),
    .A1(net389),
    .A2(net329));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_156_  (.A1(\u_ppwm/u_pwm/_077_ ),
    .A2(net330),
    .Y(\u_ppwm/u_pwm/_006_ ),
    .B1(\u_ppwm/u_pwm/_094_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_157_  (.B1(net424),
    .Y(\u_ppwm/u_pwm/_095_ ),
    .A1(net387),
    .A2(net328));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_158_  (.A1(\u_ppwm/u_pwm/_076_ ),
    .A2(net328),
    .Y(\u_ppwm/u_pwm/_007_ ),
    .B1(\u_ppwm/u_pwm/_095_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_159_  (.B1(net425),
    .Y(\u_ppwm/u_pwm/_096_ ),
    .A1(net386),
    .A2(net329));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_160_  (.A1(\u_ppwm/u_pwm/_075_ ),
    .A2(net330),
    .Y(\u_ppwm/u_pwm/_008_ ),
    .B1(\u_ppwm/u_pwm/_096_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_161_  (.B1(net425),
    .Y(\u_ppwm/u_pwm/_097_ ),
    .A1(\u_ppwm/pwm_value[9] ),
    .A2(net329));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_162_  (.A1(\u_ppwm/u_pwm/_074_ ),
    .A2(net330),
    .Y(\u_ppwm/u_pwm/_009_ ),
    .B1(\u_ppwm/u_pwm/_097_ ));
 sg13g2_and2_1 \u_ppwm/u_pwm/_163_  (.A(net625),
    .B(net630),
    .X(\u_ppwm/u_pwm/_098_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_164_  (.B1(net422),
    .Y(\u_ppwm/u_pwm/_099_ ),
    .A1(net625),
    .A2(net630));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_165_  (.A(\u_ppwm/u_pwm/_098_ ),
    .B(\u_ppwm/u_pwm/_099_ ),
    .Y(\u_ppwm/u_pwm/_010_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_166_  (.B1(net422),
    .Y(\u_ppwm/u_pwm/_100_ ),
    .A1(net535),
    .A2(\u_ppwm/u_pwm/_098_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_167_  (.A1(net535),
    .A2(\u_ppwm/u_pwm/_098_ ),
    .Y(\u_ppwm/u_pwm/_011_ ),
    .B1(\u_ppwm/u_pwm/_100_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_168_  (.A1(net535),
    .A2(\u_ppwm/u_pwm/_098_ ),
    .Y(\u_ppwm/u_pwm/_101_ ),
    .B1(net611));
 sg13g2_and4_1 \u_ppwm/u_pwm/_169_  (.A(net625),
    .B(net611),
    .C(net535),
    .D(net630),
    .X(\u_ppwm/u_pwm/_022_ ));
 sg13g2_nor3_1 \u_ppwm/u_pwm/_170_  (.A(\u_ppwm/u_pwm/_084_ ),
    .B(net612),
    .C(\u_ppwm/u_pwm/_022_ ),
    .Y(\u_ppwm/u_pwm/_012_ ));
 sg13g2_xnor2_1 \u_ppwm/u_pwm/_171_  (.Y(\u_ppwm/u_pwm/_023_ ),
    .A(net337),
    .B(\u_ppwm/u_pwm/_022_ ));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_172_  (.A(\u_ppwm/u_pwm/_084_ ),
    .B(\u_ppwm/u_pwm/_023_ ),
    .Y(\u_ppwm/u_pwm/_013_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_173_  (.A1(net337),
    .A2(\u_ppwm/u_pwm/_022_ ),
    .Y(\u_ppwm/u_pwm/_024_ ),
    .B1(net621));
 sg13g2_and3_1 \u_ppwm/u_pwm/_174_  (.X(\u_ppwm/u_pwm/_025_ ),
    .A(net621),
    .B(net337),
    .C(\u_ppwm/u_pwm/_022_ ));
 sg13g2_nor3_1 \u_ppwm/u_pwm/_175_  (.A(\u_ppwm/u_pwm/_084_ ),
    .B(net622),
    .C(\u_ppwm/u_pwm/_025_ ),
    .Y(\u_ppwm/u_pwm/_014_ ));
 sg13g2_and4_1 \u_ppwm/u_pwm/_176_  (.A(net643),
    .B(net621),
    .C(net660),
    .D(\u_ppwm/u_pwm/_022_ ),
    .X(\u_ppwm/u_pwm/_026_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_177_  (.B1(net422),
    .Y(\u_ppwm/u_pwm/_027_ ),
    .A1(net643),
    .A2(\u_ppwm/u_pwm/_025_ ));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_178_  (.A(\u_ppwm/u_pwm/_026_ ),
    .B(net644),
    .Y(\u_ppwm/u_pwm/_015_ ));
 sg13g2_or2_1 \u_ppwm/u_pwm/_179_  (.X(\u_ppwm/u_pwm/_028_ ),
    .B(\u_ppwm/u_pwm/_026_ ),
    .A(net626));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_180_  (.Y(\u_ppwm/u_pwm/_029_ ),
    .A(net626),
    .B(\u_ppwm/u_pwm/_026_ ));
 sg13g2_and3_1 \u_ppwm/u_pwm/_181_  (.X(\u_ppwm/u_pwm/_016_ ),
    .A(net422),
    .B(\u_ppwm/u_pwm/_028_ ),
    .C(\u_ppwm/u_pwm/_029_ ));
 sg13g2_nand3_1 \u_ppwm/u_pwm/_182_  (.B(net626),
    .C(\u_ppwm/u_pwm/_026_ ),
    .A(net580),
    .Y(\u_ppwm/u_pwm/_030_ ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_183_  (.Y(\u_ppwm/u_pwm/_031_ ),
    .A(net422),
    .B(\u_ppwm/u_pwm/_030_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_184_  (.A1(\u_ppwm/u_pwm/_071_ ),
    .A2(\u_ppwm/u_pwm/_029_ ),
    .Y(\u_ppwm/u_pwm/_017_ ),
    .B1(\u_ppwm/u_pwm/_031_ ));
 sg13g2_or2_1 \u_ppwm/u_pwm/_185_  (.X(\u_ppwm/u_pwm/_032_ ),
    .B(\u_ppwm/u_pwm/_030_ ),
    .A(\u_ppwm/u_pwm/_070_ ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_186_  (.Y(\u_ppwm/u_pwm/_033_ ),
    .A(net424),
    .B(\u_ppwm/u_pwm/_032_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_187_  (.A1(\u_ppwm/u_pwm/_070_ ),
    .A2(\u_ppwm/u_pwm/_030_ ),
    .Y(\u_ppwm/u_pwm/_018_ ),
    .B1(\u_ppwm/u_pwm/_033_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_188_  (.B1(net424),
    .Y(\u_ppwm/u_pwm/_034_ ),
    .A1(\u_ppwm/u_pwm/_069_ ),
    .A2(\u_ppwm/u_pwm/_032_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_189_  (.A1(\u_ppwm/u_pwm/_069_ ),
    .A2(\u_ppwm/u_pwm/_032_ ),
    .Y(\u_ppwm/u_pwm/_019_ ),
    .B1(\u_ppwm/u_pwm/_034_ ));
 sg13g2_nand3_1 \u_ppwm/u_pwm/_190_  (.B(\u_ppwm/u_pwm/counter[0] ),
    .C(net422),
    .A(net535),
    .Y(\u_ppwm/u_pwm/_035_ ));
 sg13g2_nand4_1 \u_ppwm/u_pwm/_191_  (.B(\u_ppwm/u_pwm/counter[8] ),
    .C(\u_ppwm/u_pwm/counter[5] ),
    .A(net594),
    .Y(\u_ppwm/u_pwm/_036_ ),
    .D(\u_ppwm/u_pwm/counter[4] ));
 sg13g2_nand4_1 \u_ppwm/u_pwm/_192_  (.B(\u_ppwm/u_pwm/counter[6] ),
    .C(net337),
    .A(net580),
    .Y(\u_ppwm/u_pwm/_037_ ),
    .D(\u_ppwm/u_pwm/counter[2] ));
 sg13g2_nor3_1 \u_ppwm/u_pwm/_193_  (.A(\u_ppwm/u_pwm/_035_ ),
    .B(net595),
    .C(\u_ppwm/u_pwm/_037_ ),
    .Y(\u_ppwm/u_pwm/_020_ ));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_194_  (.Y(\u_ppwm/u_pwm/_038_ ),
    .B(\u_ppwm/u_pwm/counter[2] ),
    .A_N(\u_ppwm/u_pwm/cmp_value[2] ));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_195_  (.A(\u_ppwm/u_pwm/cmp_value[3] ),
    .B_N(net337),
    .Y(\u_ppwm/u_pwm/_039_ ));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_196_  (.Y(\u_ppwm/u_pwm/_040_ ),
    .B(net337),
    .A_N(\u_ppwm/u_pwm/cmp_value[3] ));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_197_  (.A(net337),
    .B_N(\u_ppwm/u_pwm/cmp_value[3] ),
    .Y(\u_ppwm/u_pwm/_041_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_198_  (.A1(\u_ppwm/u_pwm/_038_ ),
    .A2(\u_ppwm/u_pwm/_040_ ),
    .Y(\u_ppwm/u_pwm/_042_ ),
    .B1(\u_ppwm/u_pwm/_041_ ));
 sg13g2_a221oi_1 \u_ppwm/u_pwm/_199_  (.B2(\u_ppwm/u_pwm/_073_ ),
    .C1(\u_ppwm/u_pwm/_041_ ),
    .B1(\u_ppwm/u_pwm/cmp_value[1] ),
    .A1(\u_ppwm/u_pwm/_072_ ),
    .Y(\u_ppwm/u_pwm/_043_ ),
    .A2(\u_ppwm/u_pwm/cmp_value[2] ));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_200_  (.Y(\u_ppwm/u_pwm/_044_ ),
    .B(\u_ppwm/u_pwm/counter[1] ),
    .A_N(\u_ppwm/u_pwm/cmp_value[1] ));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_201_  (.A(\u_ppwm/u_pwm/counter[0] ),
    .B_N(\u_ppwm/u_pwm/cmp_value[0] ),
    .Y(\u_ppwm/u_pwm/_045_ ));
 sg13g2_a221oi_1 \u_ppwm/u_pwm/_202_  (.B2(\u_ppwm/u_pwm/_045_ ),
    .C1(\u_ppwm/u_pwm/_039_ ),
    .B1(\u_ppwm/u_pwm/_044_ ),
    .A1(\u_ppwm/u_pwm/counter[2] ),
    .Y(\u_ppwm/u_pwm/_046_ ),
    .A2(\u_ppwm/u_pwm/_081_ ));
 sg13g2_a21o_1 \u_ppwm/u_pwm/_203_  (.A2(\u_ppwm/u_pwm/_046_ ),
    .A1(\u_ppwm/u_pwm/_043_ ),
    .B1(\u_ppwm/u_pwm/_042_ ),
    .X(\u_ppwm/u_pwm/_047_ ));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_204_  (.Y(\u_ppwm/u_pwm/_048_ ),
    .B(\u_ppwm/u_pwm/counter[7] ),
    .A_N(\u_ppwm/u_pwm/cmp_value[7] ));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_205_  (.Y(\u_ppwm/u_pwm/_049_ ),
    .B(\u_ppwm/u_pwm/counter[6] ),
    .A_N(\u_ppwm/u_pwm/cmp_value[6] ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_206_  (.Y(\u_ppwm/u_pwm/_050_ ),
    .A(\u_ppwm/u_pwm/_048_ ),
    .B(\u_ppwm/u_pwm/_049_ ));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_207_  (.Y(\u_ppwm/u_pwm/_051_ ),
    .B(\u_ppwm/u_pwm/cmp_value[7] ),
    .A_N(\u_ppwm/u_pwm/counter[7] ));
 sg13g2_nand2b_1 \u_ppwm/u_pwm/_208_  (.Y(\u_ppwm/u_pwm/_052_ ),
    .B(\u_ppwm/u_pwm/cmp_value[6] ),
    .A_N(\u_ppwm/u_pwm/counter[6] ));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_209_  (.A(\u_ppwm/u_pwm/counter[5] ),
    .B(\u_ppwm/u_pwm/_078_ ),
    .Y(\u_ppwm/u_pwm/_053_ ));
 sg13g2_nand4_1 \u_ppwm/u_pwm/_210_  (.B(\u_ppwm/u_pwm/_049_ ),
    .C(\u_ppwm/u_pwm/_051_ ),
    .A(\u_ppwm/u_pwm/_048_ ),
    .Y(\u_ppwm/u_pwm/_054_ ),
    .D(\u_ppwm/u_pwm/_052_ ));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_211_  (.A(\u_ppwm/u_pwm/_053_ ),
    .B(\u_ppwm/u_pwm/_054_ ),
    .Y(\u_ppwm/u_pwm/_055_ ));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_212_  (.A(\u_ppwm/u_pwm/cmp_value[5] ),
    .B_N(\u_ppwm/u_pwm/counter[5] ),
    .Y(\u_ppwm/u_pwm/_056_ ));
 sg13g2_a21o_1 \u_ppwm/u_pwm/_213_  (.A2(\u_ppwm/u_pwm/_079_ ),
    .A1(\u_ppwm/u_pwm/counter[4] ),
    .B1(\u_ppwm/u_pwm/_056_ ),
    .X(\u_ppwm/u_pwm/_057_ ));
 sg13g2_nor2_1 \u_ppwm/u_pwm/_214_  (.A(\u_ppwm/u_pwm/counter[4] ),
    .B(\u_ppwm/u_pwm/_079_ ),
    .Y(\u_ppwm/u_pwm/_058_ ));
 sg13g2_nor4_1 \u_ppwm/u_pwm/_215_  (.A(\u_ppwm/u_pwm/_053_ ),
    .B(\u_ppwm/u_pwm/_054_ ),
    .C(\u_ppwm/u_pwm/_057_ ),
    .D(\u_ppwm/u_pwm/_058_ ),
    .Y(\u_ppwm/u_pwm/_059_ ));
 sg13g2_and2_1 \u_ppwm/u_pwm/_216_  (.A(\u_ppwm/u_pwm/_050_ ),
    .B(\u_ppwm/u_pwm/_051_ ),
    .X(\u_ppwm/u_pwm/_060_ ));
 sg13g2_a221oi_1 \u_ppwm/u_pwm/_217_  (.B2(\u_ppwm/u_pwm/_047_ ),
    .C1(\u_ppwm/u_pwm/_060_ ),
    .B1(\u_ppwm/u_pwm/_059_ ),
    .A1(\u_ppwm/u_pwm/_055_ ),
    .Y(\u_ppwm/u_pwm/_061_ ),
    .A2(\u_ppwm/u_pwm/_057_ ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_218_  (.Y(\u_ppwm/u_pwm/_062_ ),
    .A(net604),
    .B(\u_ppwm/u_pwm/_075_ ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_219_  (.Y(\u_ppwm/u_pwm/_063_ ),
    .A(\u_ppwm/u_pwm/_069_ ),
    .B(net568));
 sg13g2_a22oi_1 \u_ppwm/u_pwm/_220_  (.Y(\u_ppwm/u_pwm/_064_ ),
    .B1(net264),
    .B2(\u_ppwm/u_pwm/_070_ ),
    .A2(net568),
    .A1(\u_ppwm/u_pwm/_069_ ));
 sg13g2_nand2_1 \u_ppwm/u_pwm/_221_  (.Y(\u_ppwm/u_pwm/_065_ ),
    .A(\u_ppwm/u_pwm/_062_ ),
    .B(\u_ppwm/u_pwm/_064_ ));
 sg13g2_nor2b_1 \u_ppwm/u_pwm/_222_  (.A(\u_ppwm/u_pwm/_062_ ),
    .B_N(\u_ppwm/u_pwm/_063_ ),
    .Y(\u_ppwm/u_pwm/_066_ ));
 sg13g2_a21oi_1 \u_ppwm/u_pwm/_223_  (.A1(net594),
    .A2(\u_ppwm/u_pwm/_074_ ),
    .Y(\u_ppwm/u_pwm/_067_ ),
    .B1(\u_ppwm/u_pwm/_066_ ));
 sg13g2_o21ai_1 \u_ppwm/u_pwm/_224_  (.B1(\u_ppwm/u_pwm/_067_ ),
    .Y(\u_ppwm/u_pwm/_068_ ),
    .A1(\u_ppwm/u_pwm/_061_ ),
    .A2(\u_ppwm/u_pwm/_065_ ));
 sg13g2_and2_1 \u_ppwm/u_pwm/_225_  (.A(net422),
    .B(\u_ppwm/u_pwm/_068_ ),
    .X(\u_ppwm/u_pwm/_021_ ));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_226_  (.RESET_B(net190),
    .D(net201),
    .Q(\u_ppwm/u_pwm/cmp_value[0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_227_  (.RESET_B(net187),
    .D(net219),
    .Q(\u_ppwm/u_pwm/cmp_value[1] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_228_  (.RESET_B(net185),
    .D(net563),
    .Q(\u_ppwm/u_pwm/cmp_value[2] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_229_  (.RESET_B(net183),
    .D(net497),
    .Q(\u_ppwm/u_pwm/cmp_value[3] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_230_  (.RESET_B(net181),
    .D(net305),
    .Q(\u_ppwm/u_pwm/cmp_value[4] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_231_  (.RESET_B(net179),
    .D(net223),
    .Q(\u_ppwm/u_pwm/cmp_value[5] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_232_  (.RESET_B(net177),
    .D(net221),
    .Q(\u_ppwm/u_pwm/cmp_value[6] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_233_  (.RESET_B(net197),
    .D(net250),
    .Q(\u_ppwm/u_pwm/cmp_value[7] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_234_  (.RESET_B(net195),
    .D(net265),
    .Q(\u_ppwm/u_pwm/cmp_value[8] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_235_  (.RESET_B(net193),
    .D(net569),
    .Q(\u_ppwm/u_pwm/cmp_value[9] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_236_  (.RESET_B(net191),
    .D(\u_ppwm/u_pwm/_010_ ),
    .Q(\u_ppwm/u_pwm/counter[0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_237_  (.RESET_B(net189),
    .D(net536),
    .Q(\u_ppwm/u_pwm/counter[1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_238_  (.RESET_B(net186),
    .D(net613),
    .Q(\u_ppwm/u_pwm/counter[2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_239_  (.RESET_B(net182),
    .D(\u_ppwm/u_pwm/_013_ ),
    .Q(\u_ppwm/u_pwm/counter[3] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_240_  (.RESET_B(net178),
    .D(net623),
    .Q(\u_ppwm/u_pwm/counter[4] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_241_  (.RESET_B(net196),
    .D(net645),
    .Q(\u_ppwm/u_pwm/counter[5] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_242_  (.RESET_B(net192),
    .D(\u_ppwm/u_pwm/_016_ ),
    .Q(\u_ppwm/u_pwm/counter[6] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_243_  (.RESET_B(net188),
    .D(net581),
    .Q(\u_ppwm/u_pwm/counter[7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_244_  (.RESET_B(net180),
    .D(net605),
    .Q(\u_ppwm/u_pwm/counter[8] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_245_  (.RESET_B(net194),
    .D(\u_ppwm/u_pwm/_019_ ),
    .Q(\u_ppwm/u_pwm/counter[9] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 \u_ppwm/u_pwm/_246_  (.RESET_B(net184),
    .D(net596),
    .Q(\u_ppwm/period_start ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 \u_ppwm/u_pwm/_247_  (.RESET_B(net176),
    .D(\u_ppwm/u_pwm/_021_ ),
    .Q(net2),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_tiehi \u_ppwm/u_pwm/_232__177  (.L_HI(net177));
 sg13g2_tiehi \u_ppwm/u_pwm/_240__178  (.L_HI(net178));
 sg13g2_tiehi \u_ppwm/u_pwm/_231__179  (.L_HI(net179));
 sg13g2_tiehi \u_ppwm/u_pwm/_244__180  (.L_HI(net180));
 sg13g2_tiehi \u_ppwm/u_pwm/_230__181  (.L_HI(net181));
 sg13g2_tiehi \u_ppwm/u_pwm/_239__182  (.L_HI(net182));
 sg13g2_tiehi \u_ppwm/u_pwm/_229__183  (.L_HI(net183));
 sg13g2_tiehi \u_ppwm/u_pwm/_246__184  (.L_HI(net184));
 sg13g2_tiehi \u_ppwm/u_pwm/_228__185  (.L_HI(net185));
 sg13g2_tiehi \u_ppwm/u_pwm/_238__186  (.L_HI(net186));
 sg13g2_tiehi \u_ppwm/u_pwm/_227__187  (.L_HI(net187));
 sg13g2_tiehi \u_ppwm/u_pwm/_243__188  (.L_HI(net188));
 sg13g2_tiehi \u_ppwm/u_pwm/_237__189  (.L_HI(net189));
 sg13g2_tiehi \u_ppwm/u_pwm/_226__190  (.L_HI(net190));
 sg13g2_tiehi \u_ppwm/u_pwm/_236__191  (.L_HI(net191));
 sg13g2_tiehi \u_ppwm/u_pwm/_242__192  (.L_HI(net192));
 sg13g2_tiehi \u_ppwm/u_pwm/_235__193  (.L_HI(net193));
 sg13g2_tiehi \u_ppwm/u_pwm/_245__194  (.L_HI(net194));
 sg13g2_tiehi \u_ppwm/u_pwm/_234__195  (.L_HI(net195));
 sg13g2_tiehi \u_ppwm/u_pwm/_241__196  (.L_HI(net196));
 sg13g2_tiehi \u_ppwm/u_pwm/_233__197  (.L_HI(net197));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 fanout307 (.A(\u_ppwm/u_ex/_294_ ),
    .X(net307));
 sg13g2_buf_1 fanout308 (.A(\u_ppwm/u_ex/_294_ ),
    .X(net308));
 sg13g2_buf_8 fanout309 (.A(\u_ppwm/u_ex/_214_ ),
    .X(net309));
 sg13g2_buf_8 fanout310 (.A(\u_ppwm/u_ex/_213_ ),
    .X(net310));
 sg13g2_buf_8 fanout311 (.A(net312),
    .X(net311));
 sg13g2_buf_8 fanout312 (.A(\u_ppwm/u_ex/_227_ ),
    .X(net312));
 sg13g2_buf_8 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_8 fanout314 (.A(\u_ppwm/u_ex/_221_ ),
    .X(net314));
 sg13g2_buf_8 fanout315 (.A(\u_ppwm/u_ex/_217_ ),
    .X(net315));
 sg13g2_buf_8 fanout316 (.A(\u_ppwm/u_ex/_216_ ),
    .X(net316));
 sg13g2_buf_8 fanout317 (.A(\u_ppwm/u_ex/_215_ ),
    .X(net317));
 sg13g2_buf_8 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_8 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_8 fanout320 (.A(\u_ppwm/instr[6] ),
    .X(net320));
 sg13g2_buf_8 fanout321 (.A(net322),
    .X(net321));
 sg13g2_buf_8 fanout322 (.A(\u_ppwm/instr[6] ),
    .X(net322));
 sg13g2_buf_8 fanout323 (.A(\u_ppwm/instr[5] ),
    .X(net323));
 sg13g2_buf_1 fanout324 (.A(\u_ppwm/instr[5] ),
    .X(net324));
 sg13g2_buf_8 fanout325 (.A(net326),
    .X(net325));
 sg13g2_buf_8 fanout326 (.A(\u_ppwm/instr[4] ),
    .X(net326));
 sg13g2_buf_8 fanout327 (.A(\u_ppwm/instr[3] ),
    .X(net327));
 sg13g2_buf_8 fanout328 (.A(\u_ppwm/u_pwm/_087_ ),
    .X(net328));
 sg13g2_buf_1 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_8 fanout330 (.A(\u_ppwm/u_pwm/_087_ ),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(\u_ppwm/u_global_counter/_041_ ),
    .X(net331));
 sg13g2_buf_8 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_8 fanout333 (.A(\u_ppwm/u_mem/_0241_ ),
    .X(net333));
 sg13g2_buf_8 fanout334 (.A(net335),
    .X(net334));
 sg13g2_buf_8 fanout335 (.A(\u_ppwm/u_mem/_0240_ ),
    .X(net335));
 sg13g2_buf_8 fanout336 (.A(net661),
    .X(net336));
 sg13g2_buf_8 fanout337 (.A(net660),
    .X(net337));
 sg13g2_buf_8 fanout338 (.A(net343),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(net343),
    .X(net339));
 sg13g2_buf_8 fanout340 (.A(net342),
    .X(net340));
 sg13g2_buf_1 fanout341 (.A(net342),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_8 fanout343 (.A(net376),
    .X(net343));
 sg13g2_buf_8 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_8 fanout345 (.A(net376),
    .X(net345));
 sg13g2_buf_8 fanout346 (.A(net347),
    .X(net346));
 sg13g2_buf_8 fanout347 (.A(net357),
    .X(net347));
 sg13g2_buf_8 fanout348 (.A(net352),
    .X(net348));
 sg13g2_buf_1 fanout349 (.A(net352),
    .X(net349));
 sg13g2_buf_8 fanout350 (.A(net352),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(net357),
    .X(net352));
 sg13g2_buf_8 fanout353 (.A(net357),
    .X(net353));
 sg13g2_buf_1 fanout354 (.A(net357),
    .X(net354));
 sg13g2_buf_8 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_8 fanout356 (.A(net357),
    .X(net356));
 sg13g2_buf_8 fanout357 (.A(net376),
    .X(net357));
 sg13g2_buf_8 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_1 fanout359 (.A(net376),
    .X(net359));
 sg13g2_buf_8 fanout360 (.A(net363),
    .X(net360));
 sg13g2_buf_1 fanout361 (.A(net363),
    .X(net361));
 sg13g2_buf_8 fanout362 (.A(net363),
    .X(net362));
 sg13g2_buf_8 fanout363 (.A(net376),
    .X(net363));
 sg13g2_buf_8 fanout364 (.A(net375),
    .X(net364));
 sg13g2_buf_1 fanout365 (.A(net375),
    .X(net365));
 sg13g2_buf_8 fanout366 (.A(net369),
    .X(net366));
 sg13g2_buf_1 fanout367 (.A(net369),
    .X(net367));
 sg13g2_buf_8 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_8 fanout369 (.A(net375),
    .X(net369));
 sg13g2_buf_8 fanout370 (.A(net371),
    .X(net370));
 sg13g2_buf_8 fanout371 (.A(net372),
    .X(net371));
 sg13g2_buf_8 fanout372 (.A(net375),
    .X(net372));
 sg13g2_buf_8 fanout373 (.A(net374),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_8 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_8 fanout376 (.A(\u_ppwm/u_mem/state_q[2] ),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(net631),
    .X(net377));
 sg13g2_buf_8 fanout378 (.A(net648),
    .X(net378));
 sg13g2_buf_8 fanout379 (.A(net646),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(net639),
    .X(net380));
 sg13g2_buf_8 fanout381 (.A(net663),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(net636),
    .X(net382));
 sg13g2_buf_8 fanout383 (.A(\u_ppwm/u_ex/reg_value_q[3] ),
    .X(net383));
 sg13g2_buf_8 fanout384 (.A(net658),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(net671),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(net676),
    .X(net386));
 sg13g2_buf_8 fanout387 (.A(net673),
    .X(net387));
 sg13g2_buf_1 fanout388 (.A(\u_ppwm/pwm_value[7] ),
    .X(net388));
 sg13g2_buf_8 fanout389 (.A(net668),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(\u_ppwm/pwm_value[6] ),
    .X(net390));
 sg13g2_buf_8 fanout391 (.A(net675),
    .X(net391));
 sg13g2_buf_8 fanout392 (.A(net666),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(\u_ppwm/pwm_value[4] ),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(net664),
    .X(net394));
 sg13g2_buf_1 fanout395 (.A(\u_ppwm/pwm_value[3] ),
    .X(net395));
 sg13g2_buf_8 fanout396 (.A(net662),
    .X(net396));
 sg13g2_buf_1 fanout397 (.A(\u_ppwm/pwm_value[2] ),
    .X(net397));
 sg13g2_buf_8 fanout398 (.A(net670),
    .X(net398));
 sg13g2_buf_1 fanout399 (.A(\u_ppwm/pwm_value[1] ),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(\u_ppwm/pc[3] ),
    .X(net400));
 sg13g2_buf_1 fanout401 (.A(\u_ppwm/pc[3] ),
    .X(net401));
 sg13g2_buf_8 fanout402 (.A(net638),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(\u_ppwm/pc[2] ),
    .X(net403));
 sg13g2_buf_8 fanout404 (.A(net406),
    .X(net404));
 sg13g2_buf_1 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_8 fanout406 (.A(net409),
    .X(net406));
 sg13g2_buf_8 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_8 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(\u_ppwm/pc[1] ),
    .X(net409));
 sg13g2_buf_8 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_8 fanout411 (.A(net414),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(net413),
    .X(net412));
 sg13g2_buf_8 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_8 fanout414 (.A(net421),
    .X(net414));
 sg13g2_buf_8 fanout415 (.A(net421),
    .X(net415));
 sg13g2_buf_8 fanout416 (.A(net421),
    .X(net416));
 sg13g2_buf_8 fanout417 (.A(net420),
    .X(net417));
 sg13g2_buf_8 fanout418 (.A(net420),
    .X(net418));
 sg13g2_buf_1 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(net421),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(net672),
    .X(net421));
 sg13g2_buf_8 fanout422 (.A(net437),
    .X(net422));
 sg13g2_buf_8 fanout423 (.A(net437),
    .X(net423));
 sg13g2_buf_8 fanout424 (.A(net427),
    .X(net424));
 sg13g2_buf_1 fanout425 (.A(net427),
    .X(net425));
 sg13g2_buf_8 fanout426 (.A(net427),
    .X(net426));
 sg13g2_buf_8 fanout427 (.A(net437),
    .X(net427));
 sg13g2_buf_8 fanout428 (.A(net432),
    .X(net428));
 sg13g2_buf_8 fanout429 (.A(net432),
    .X(net429));
 sg13g2_buf_8 fanout430 (.A(net431),
    .X(net430));
 sg13g2_buf_8 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_8 fanout432 (.A(net436),
    .X(net432));
 sg13g2_buf_8 fanout433 (.A(net436),
    .X(net433));
 sg13g2_buf_8 fanout434 (.A(net435),
    .X(net434));
 sg13g2_buf_8 fanout435 (.A(net436),
    .X(net435));
 sg13g2_buf_8 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_8 fanout437 (.A(net452),
    .X(net437));
 sg13g2_buf_8 fanout438 (.A(net439),
    .X(net438));
 sg13g2_buf_8 fanout439 (.A(net442),
    .X(net439));
 sg13g2_buf_8 fanout440 (.A(net442),
    .X(net440));
 sg13g2_buf_8 fanout441 (.A(net442),
    .X(net441));
 sg13g2_buf_8 fanout442 (.A(net452),
    .X(net442));
 sg13g2_buf_8 fanout443 (.A(net446),
    .X(net443));
 sg13g2_buf_8 fanout444 (.A(net445),
    .X(net444));
 sg13g2_buf_8 fanout445 (.A(net446),
    .X(net445));
 sg13g2_buf_8 fanout446 (.A(net452),
    .X(net446));
 sg13g2_buf_8 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_8 fanout448 (.A(net451),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(net451),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(net451),
    .X(net450));
 sg13g2_buf_8 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_8 fanout452 (.A(rst_n),
    .X(net452));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_tielo heichips25_ppwm_3 (.L_LO(net3));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_5_26__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_ppwm/global_counter_high[16] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_ppwm/u_global_counter/_016_ ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_ppwm/u_pwm/cmp_value[0] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold4 (.A(\u_ppwm/u_pwm/_000_ ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_ppwm/global_counter_high[6] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_ppwm/u_global_counter/_006_ ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold7 (.A(\u_ppwm/global_counter_high[19] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold8 (.A(\u_ppwm/u_global_counter/_019_ ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_ppwm/u_mem/_0003_ ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_ppwm/u_mem/_0117_ ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_ppwm/u_mem/memory[68] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_ppwm/u_mem/_0074_ ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_ppwm/u_mem/memory[90] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_ppwm/u_mem/_0096_ ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_ppwm/u_mem/memory[99] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_ppwm/u_mem/_0105_ ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold17 (.A(\u_ppwm/u_mem/memory[57] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_ppwm/u_mem/_0063_ ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_ppwm/u_mem/memory[32] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold20 (.A(\u_ppwm/u_mem/_0038_ ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_ppwm/u_pwm/cmp_value[1] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold22 (.A(\u_ppwm/u_pwm/_001_ ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_ppwm/u_pwm/cmp_value[6] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_ppwm/u_pwm/_006_ ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_ppwm/u_pwm/cmp_value[5] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold26 (.A(\u_ppwm/u_pwm/_005_ ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_ppwm/u_mem/memory[58] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold28 (.A(\u_ppwm/u_mem/memory[82] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_ppwm/u_mem/_0088_ ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold30 (.A(\u_ppwm/global_counter_high[10] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_ppwm/u_global_counter/_010_ ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold32 (.A(\u_ppwm/u_mem/memory[78] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_ppwm/u_mem/_0084_ ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u_ppwm/u_mem/memory[86] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_ppwm/u_mem/_0092_ ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u_ppwm/u_mem/memory[106] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_ppwm/u_mem/_0112_ ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_ppwm/u_mem/memory[28] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u_ppwm/u_mem/_0034_ ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold40 (.A(\u_ppwm/u_mem/memory[51] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_ppwm/u_mem/_0057_ ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u_ppwm/u_mem/memory[81] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_ppwm/u_mem/_0087_ ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold44 (.A(\u_ppwm/u_mem/memory[9] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_ppwm/u_mem/_0015_ ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold46 (.A(\u_ppwm/u_mem/memory[67] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_ppwm/u_mem/_0073_ ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_ppwm/u_mem/memory[89] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_ppwm/u_mem/_0095_ ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u_ppwm/u_mem/memory[48] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_ppwm/u_mem/_0054_ ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u_ppwm/u_pwm/cmp_value[7] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_ppwm/u_pwm/_007_ ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u_ppwm/global_counter_high[2] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_ppwm/u_global_counter/_002_ ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u_ppwm/u_mem/memory[59] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u_ppwm/u_mem/memory[27] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold58 (.A(\u_ppwm/u_mem/_0033_ ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold59 (.A(\u_ppwm/u_mem/memory[54] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_ppwm/u_mem/_0060_ ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold61 (.A(\u_ppwm/u_mem/memory[88] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u_ppwm/u_mem/_0094_ ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold63 (.A(\u_ppwm/u_mem/memory[50] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_ppwm/u_mem/_0056_ ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold65 (.A(\u_ppwm/u_mem/memory[98] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_ppwm/u_mem/_0104_ ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold67 (.A(\u_ppwm/u_pwm/cmp_value[8] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_ppwm/u_pwm/_008_ ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold69 (.A(\u_ppwm/u_mem/memory[91] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold70 (.A(\u_ppwm/u_mem/_0097_ ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold71 (.A(\u_ppwm/global_counter_high[0] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold72 (.A(\u_ppwm/u_global_counter/_000_ ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold73 (.A(\u_ppwm/u_mem/memory[65] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold74 (.A(\u_ppwm/u_mem/_0071_ ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold75 (.A(\u_ppwm/u_mem/memory[33] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold76 (.A(\u_ppwm/u_mem/_0039_ ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold77 (.A(\u_ppwm/u_mem/memory[93] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_ppwm/u_mem/_0099_ ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold79 (.A(\u_ppwm/u_mem/memory[71] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_ppwm/u_mem/_0077_ ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold81 (.A(\u_ppwm/u_mem/memory[72] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_ppwm/u_mem/_0078_ ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold83 (.A(\u_ppwm/u_mem/memory[39] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_ppwm/u_mem/_0045_ ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold85 (.A(\u_ppwm/u_mem/memory[56] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_ppwm/u_mem/_0062_ ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold87 (.A(\u_ppwm/u_mem/memory[87] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_ppwm/u_mem/_0093_ ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold89 (.A(\u_ppwm/u_mem/memory[100] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold90 (.A(\u_ppwm/u_mem/memory[61] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold91 (.A(\u_ppwm/u_mem/_0067_ ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_ppwm/u_mem/memory[35] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold93 (.A(\u_ppwm/u_mem/_0041_ ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold94 (.A(\u_ppwm/global_counter_high[8] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_ppwm/u_global_counter/_008_ ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold96 (.A(\u_ppwm/u_mem/memory[74] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_ppwm/u_mem/_0080_ ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold98 (.A(\u_ppwm/u_mem/memory[95] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold99 (.A(\u_ppwm/u_mem/_0101_ ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold100 (.A(\u_ppwm/u_mem/memory[45] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold101 (.A(\u_ppwm/u_mem/_0051_ ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_ppwm/u_mem/memory[25] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold103 (.A(\u_ppwm/u_mem/_0031_ ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold104 (.A(\u_ppwm/u_mem/memory[18] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold105 (.A(\u_ppwm/u_mem/_0024_ ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold106 (.A(\u_ppwm/u_mem/memory[66] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold107 (.A(\u_ppwm/u_pwm/cmp_value[4] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold108 (.A(\u_ppwm/u_pwm/_004_ ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_ppwm/u_mem/memory[52] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold110 (.A(\u_ppwm/u_mem/memory[70] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold111 (.A(\u_ppwm/u_mem/_0076_ ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold112 (.A(\u_ppwm/u_mem/memory[47] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_ppwm/u_mem/_0053_ ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold114 (.A(\u_ppwm/u_mem/memory[46] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold115 (.A(\u_ppwm/u_mem/memory[94] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold116 (.A(\u_ppwm/u_mem/memory[37] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold117 (.A(\u_ppwm/u_mem/_0043_ ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold118 (.A(\u_ppwm/global_counter_high[7] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold119 (.A(\u_ppwm/u_global_counter/_036_ ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold120 (.A(\u_ppwm/u_global_counter/_007_ ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold121 (.A(\u_ppwm/u_mem/memory[11] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold122 (.A(\u_ppwm/u_mem/_0017_ ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_ppwm/u_mem/memory[38] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold124 (.A(\u_ppwm/u_mem/memory[64] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold125 (.A(\u_ppwm/u_mem/_0070_ ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold126 (.A(\u_ppwm/u_mem/memory[12] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_ppwm/u_mem/_0018_ ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_ppwm/u_mem/memory[102] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold129 (.A(\u_ppwm/u_mem/_0108_ ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_ppwm/u_mem/memory[96] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold131 (.A(\u_ppwm/u_mem/_0102_ ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_ppwm/u_mem/memory[24] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold133 (.A(\u_ppwm/u_mem/_0030_ ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold134 (.A(\u_ppwm/u_mem/memory[104] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold135 (.A(\u_ppwm/u_mem/_0110_ ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_ppwm/u_mem/memory[21] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold137 (.A(\u_ppwm/u_mem/_0027_ ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold138 (.A(\u_ppwm/u_mem/memory[7] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_ppwm/u_mem/_0013_ ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold140 (.A(\u_ppwm/u_mem/memory[17] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_ppwm/u_mem/_0023_ ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold142 (.A(\u_ppwm/u_mem/memory[85] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold143 (.A(\u_ppwm/u_mem/_0091_ ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold144 (.A(\u_ppwm/u_mem/memory[63] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_ppwm/u_mem/_0069_ ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_ppwm/u_mem/memory[97] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_ppwm/u_mem/_0103_ ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold148 (.A(\u_ppwm/u_mem/memory[13] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold149 (.A(\u_ppwm/u_mem/_0019_ ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold150 (.A(\u_ppwm/u_mem/memory[60] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold151 (.A(\u_ppwm/u_mem/memory[36] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_ppwm/u_mem/_0042_ ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_ppwm/u_pwm/cmp_value[3] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold154 (.A(\u_ppwm/u_pwm/_003_ ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_ppwm/u_mem/memory[92] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold156 (.A(\u_ppwm/u_mem/_0098_ ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_ppwm/u_mem/memory[22] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold158 (.A(\u_ppwm/u_mem/memory[3] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_ppwm/u_mem/_0009_ ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_ppwm/u_mem/memory[19] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold161 (.A(\u_ppwm/u_mem/_0025_ ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_ppwm/u_mem/memory[23] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold163 (.A(\u_ppwm/u_mem/memory[14] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold164 (.A(\u_ppwm/u_mem/_0020_ ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold165 (.A(\u_ppwm/u_mem/memory[80] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold166 (.A(\u_ppwm/u_mem/_0086_ ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold167 (.A(\u_ppwm/u_mem/memory[73] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold168 (.A(\u_ppwm/u_mem/memory[1] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_ppwm/u_mem/_0007_ ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold170 (.A(\u_ppwm/u_mem/state_q[0] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold171 (.A(\u_ppwm/u_mem/_0004_ ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold172 (.A(\u_ppwm/u_mem/memory[49] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold173 (.A(\u_ppwm/u_mem/memory[83] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold174 (.A(\u_ppwm/u_mem/memory[31] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold175 (.A(\u_ppwm/u_mem/_0037_ ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_ppwm/u_mem/memory[43] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold177 (.A(\u_ppwm/u_mem/_0049_ ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold178 (.A(\u_ppwm/u_mem/_0002_ ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_ppwm/u_mem/_0116_ ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold180 (.A(\u_ppwm/u_mem/memory[10] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_ppwm/u_mem/memory[75] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold182 (.A(\u_ppwm/u_mem/memory[77] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold183 (.A(\u_ppwm/u_mem/_0083_ ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold184 (.A(\u_ppwm/u_mem/memory[4] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold185 (.A(\u_ppwm/global_counter_high[4] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_ppwm/u_global_counter/_004_ ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold187 (.A(\u_ppwm/u_mem/memory[30] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold188 (.A(\u_ppwm/u_mem/_0036_ ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_ppwm/u_mem/memory[5] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold190 (.A(\u_ppwm/u_mem/_0011_ ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold191 (.A(\u_ppwm/u_mem/memory[103] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold192 (.A(\u_ppwm/u_pwm/counter[1] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_ppwm/u_pwm/_011_ ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold194 (.A(\u_ppwm/u_mem/memory[20] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_ppwm/u_mem/memory[79] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold196 (.A(\u_ppwm/u_mem/memory[42] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_ppwm/u_mem/_0048_ ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold198 (.A(\u_ppwm/u_mem/memory[41] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_ppwm/u_mem/_0047_ ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold200 (.A(\u_ppwm/u_mem/memory[107] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold201 (.A(\u_ppwm/u_mem/memory[76] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold202 (.A(\u_ppwm/u_mem/memory[40] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold203 (.A(\u_ppwm/global_counter_high[3] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold204 (.A(\u_ppwm/u_global_counter/_003_ ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_ppwm/u_mem/memory[44] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold206 (.A(\u_ppwm/u_mem/bit_count[6] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold207 (.A(\u_ppwm/u_mem/_0489_ ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold208 (.A(\u_ppwm/u_mem/_0125_ ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold209 (.A(\u_ppwm/global_counter_high[14] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold210 (.A(\u_ppwm/u_global_counter/_045_ ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold211 (.A(\u_ppwm/u_global_counter/_014_ ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold212 (.A(\u_ppwm/global_counter_high[12] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold213 (.A(\u_ppwm/u_global_counter/_042_ ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold214 (.A(\u_ppwm/u_global_counter/_012_ ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold215 (.A(\u_ppwm/u_mem/_0000_ ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold216 (.A(\u_ppwm/u_mem/memory[55] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold217 (.A(\u_ppwm/u_mem/memory[8] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold218 (.A(\u_ppwm/u_mem/_0014_ ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold219 (.A(\u_ppwm/u_pwm/cmp_value[2] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold220 (.A(\u_ppwm/u_pwm/_002_ ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold221 (.A(\u_ppwm/global_counter_high[18] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold222 (.A(\u_ppwm/u_global_counter/_018_ ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_ppwm/u_mem/memory[105] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold224 (.A(\u_ppwm/u_mem/_0111_ ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold225 (.A(\u_ppwm/u_pwm/cmp_value[9] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold226 (.A(\u_ppwm/u_pwm/_009_ ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold227 (.A(\u_ppwm/u_mem/memory[26] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold228 (.A(\u_ppwm/u_mem/_0032_ ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold229 (.A(\u_ppwm/u_ex/state_q[0] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold230 (.A(\u_ppwm/u_ex/_000_ ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold231 (.A(\u_ppwm/u_mem/memory[84] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_ppwm/u_mem/memory[29] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold233 (.A(\u_ppwm/u_mem/memory[53] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold234 (.A(\u_ppwm/global_counter_high[15] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold235 (.A(\u_ppwm/u_global_counter/_015_ ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold236 (.A(\u_ppwm/u_mem/memory[101] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold237 (.A(\u_ppwm/u_pwm/counter[7] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold238 (.A(\u_ppwm/u_pwm/_017_ ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold239 (.A(\u_ppwm/u_mem/bit_count[2] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold240 (.A(\u_ppwm/u_mem/_0481_ ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold241 (.A(\u_ppwm/u_mem/_0121_ ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold242 (.A(\u_ppwm/u_mem/memory[2] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold243 (.A(\u_ppwm/global_counter_high[5] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold244 (.A(\u_ppwm/u_global_counter/_033_ ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold245 (.A(\u_ppwm/u_global_counter/_005_ ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold246 (.A(\u_ppwm/u_mem/memory[15] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold247 (.A(\u_ppwm/u_mem/_0021_ ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold248 (.A(\u_ppwm/u_mem/memory[16] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold249 (.A(\u_ppwm/u_mem/_0001_ ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold250 (.A(\u_ppwm/u_mem/_0115_ ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold251 (.A(\u_ppwm/u_pwm/counter[9] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold252 (.A(\u_ppwm/u_pwm/_036_ ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold253 (.A(\u_ppwm/u_pwm/_020_ ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold254 (.A(\u_ppwm/u_mem/bit_count[5] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold255 (.A(\u_ppwm/u_mem/_0487_ ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold256 (.A(\u_ppwm/u_mem/_0124_ ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold257 (.A(\u_ppwm/u_mem/memory[6] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold258 (.A(\u_ppwm/u_mem/_0012_ ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold259 (.A(\u_ppwm/u_mem/bit_count[4] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold260 (.A(\u_ppwm/u_mem/_0247_ ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold261 (.A(\u_ppwm/u_pwm/counter[8] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold262 (.A(\u_ppwm/u_pwm/_018_ ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold263 (.A(\u_ppwm/u_mem/memory[34] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold264 (.A(\u_ppwm/u_ex/state_q[1] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold265 (.A(\u_ppwm/u_ex/_052_ ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold266 (.A(\u_ppwm/global_counter_high[11] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold267 (.A(\u_ppwm/u_global_counter/_011_ ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold268 (.A(\u_ppwm/u_pwm/counter[2] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold269 (.A(\u_ppwm/u_pwm/_101_ ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold270 (.A(\u_ppwm/u_pwm/_012_ ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold271 (.A(\u_ppwm/global_counter_high[17] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold272 (.A(\u_ppwm/global_counter_high[13] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold273 (.A(\u_ppwm/u_global_counter/_013_ ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold274 (.A(\u_ppwm/u_mem/memory[62] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold275 (.A(\u_ppwm/u_mem/bit_count[0] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold276 (.A(\u_ppwm/u_mem/bit_count[1] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold277 (.A(\u_ppwm/u_mem/memory[69] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold278 (.A(\u_ppwm/u_pwm/counter[4] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold279 (.A(\u_ppwm/u_pwm/_024_ ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold280 (.A(\u_ppwm/u_pwm/_014_ ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold281 (.A(\u_ppwm/u_mem/bit_count[3] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold282 (.A(\u_ppwm/mem_write_done ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold283 (.A(\u_ppwm/u_pwm/counter[6] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold284 (.A(\u_ppwm/u_ex/cmp_flag_q ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold285 (.A(\u_ppwm/u_ex/_210_ ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold286 (.A(\u_ppwm/u_ex/_007_ ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold287 (.A(\u_ppwm/u_pwm/counter[0] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold288 (.A(\u_ppwm/u_ex/state_q[2] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold289 (.A(\u_ppwm/u_ex/_084_ ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold290 (.A(\u_ppwm/u_ex/_006_ ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold291 (.A(\u_ppwm/u_ex/reg_value_q[1] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold292 (.A(\u_ppwm/u_ex/_018_ ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold293 (.A(\u_ppwm/u_ex/reg_value_q[4] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold294 (.A(\u_ppwm/u_ex/_022_ ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_ppwm/pc[2] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold296 (.A(\u_ppwm/u_ex/reg_value_q[6] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold297 (.A(\u_ppwm/u_ex/_024_ ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold298 (.A(\u_ppwm/u_ex/reg_value_q[0] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold299 (.A(\u_ppwm/u_ex/_019_ ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold300 (.A(\u_ppwm/u_pwm/counter[5] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold301 (.A(\u_ppwm/u_pwm/_027_ ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold302 (.A(\u_ppwm/u_pwm/_015_ ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold303 (.A(\u_ppwm/u_ex/reg_value_q[8] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold304 (.A(\u_ppwm/u_ex/_026_ ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold305 (.A(\u_ppwm/u_ex/reg_value_q[9] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold306 (.A(\u_ppwm/pwm_value[0] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold307 (.A(\u_ppwm/u_ex/_008_ ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold308 (.A(\u_ppwm/pwm_value[9] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold309 (.A(\u_ppwm/u_ex/_017_ ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold310 (.A(\u_ppwm/u_ex/reg_value_q[7] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold311 (.A(\u_ppwm/global_counter_high[1] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold312 (.A(\u_ppwm/u_global_counter/_028_ ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold313 (.A(\u_ppwm/u_global_counter/_001_ ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold314 (.A(\u_ppwm/global_counter_high[9] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold315 (.A(\u_ppwm/u_ex/reg_value_q[2] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold316 (.A(\u_ppwm/u_ex/_021_ ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold317 (.A(\u_ppwm/u_pwm/counter[3] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold318 (.A(\u_ppwm/period_start ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold319 (.A(\u_ppwm/pwm_value[2] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold320 (.A(\u_ppwm/u_ex/reg_value_q[5] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold321 (.A(\u_ppwm/pwm_value[3] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold322 (.A(\u_ppwm/u_ex/_011_ ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold323 (.A(\u_ppwm/pwm_value[4] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold324 (.A(\u_ppwm/u_ex/_012_ ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold325 (.A(\u_ppwm/pwm_value[6] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold326 (.A(\u_ppwm/u_ex/_014_ ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold327 (.A(\u_ppwm/pwm_value[1] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold328 (.A(\u_ppwm/u_ex/reg_value_q[1] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold329 (.A(\u_ppwm/pc[0] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold330 (.A(\u_ppwm/pwm_value[7] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold331 (.A(\u_ppwm/u_ex/_015_ ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold332 (.A(\u_ppwm/pwm_value[5] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold333 (.A(\u_ppwm/pwm_value[8] ),
    .X(net676));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_fill_1 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_fill_1 FILLER_0_109 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_fill_1 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_8 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_fill_2 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_414 ();
 sg13g2_decap_8 FILLER_0_421 ();
 sg13g2_decap_8 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_0_435 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_decap_8 FILLER_0_449 ();
 sg13g2_decap_8 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_463 ();
 sg13g2_decap_8 FILLER_0_470 ();
 sg13g2_decap_8 FILLER_0_477 ();
 sg13g2_decap_8 FILLER_0_484 ();
 sg13g2_decap_8 FILLER_0_491 ();
 sg13g2_decap_8 FILLER_0_498 ();
 sg13g2_decap_8 FILLER_0_505 ();
 sg13g2_decap_8 FILLER_0_512 ();
 sg13g2_decap_8 FILLER_0_519 ();
 sg13g2_decap_8 FILLER_0_526 ();
 sg13g2_decap_8 FILLER_0_533 ();
 sg13g2_decap_8 FILLER_0_540 ();
 sg13g2_decap_8 FILLER_0_547 ();
 sg13g2_decap_8 FILLER_0_554 ();
 sg13g2_decap_8 FILLER_0_561 ();
 sg13g2_decap_8 FILLER_0_568 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_decap_8 FILLER_0_582 ();
 sg13g2_decap_8 FILLER_0_589 ();
 sg13g2_decap_8 FILLER_0_596 ();
 sg13g2_decap_8 FILLER_0_603 ();
 sg13g2_decap_8 FILLER_0_610 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_decap_8 FILLER_0_624 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_decap_8 FILLER_0_638 ();
 sg13g2_decap_8 FILLER_0_645 ();
 sg13g2_decap_8 FILLER_0_652 ();
 sg13g2_decap_8 FILLER_0_659 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_decap_8 FILLER_0_680 ();
 sg13g2_decap_8 FILLER_0_687 ();
 sg13g2_decap_8 FILLER_0_694 ();
 sg13g2_decap_8 FILLER_0_701 ();
 sg13g2_decap_8 FILLER_0_708 ();
 sg13g2_decap_8 FILLER_0_715 ();
 sg13g2_decap_8 FILLER_0_722 ();
 sg13g2_decap_8 FILLER_0_729 ();
 sg13g2_decap_8 FILLER_0_736 ();
 sg13g2_decap_8 FILLER_0_743 ();
 sg13g2_decap_8 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_757 ();
 sg13g2_decap_8 FILLER_0_764 ();
 sg13g2_decap_8 FILLER_0_771 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_decap_8 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_799 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_820 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_834 ();
 sg13g2_decap_8 FILLER_0_841 ();
 sg13g2_decap_8 FILLER_0_848 ();
 sg13g2_decap_8 FILLER_0_855 ();
 sg13g2_decap_8 FILLER_0_862 ();
 sg13g2_decap_8 FILLER_0_869 ();
 sg13g2_decap_8 FILLER_0_876 ();
 sg13g2_decap_8 FILLER_0_883 ();
 sg13g2_decap_8 FILLER_0_890 ();
 sg13g2_decap_8 FILLER_0_897 ();
 sg13g2_decap_8 FILLER_0_904 ();
 sg13g2_decap_8 FILLER_0_911 ();
 sg13g2_decap_8 FILLER_0_918 ();
 sg13g2_decap_8 FILLER_0_925 ();
 sg13g2_decap_8 FILLER_0_932 ();
 sg13g2_decap_8 FILLER_0_939 ();
 sg13g2_decap_8 FILLER_0_946 ();
 sg13g2_decap_8 FILLER_0_953 ();
 sg13g2_decap_8 FILLER_0_960 ();
 sg13g2_decap_8 FILLER_0_967 ();
 sg13g2_decap_8 FILLER_0_974 ();
 sg13g2_decap_8 FILLER_0_981 ();
 sg13g2_decap_8 FILLER_0_988 ();
 sg13g2_decap_8 FILLER_0_995 ();
 sg13g2_decap_8 FILLER_0_1002 ();
 sg13g2_decap_8 FILLER_0_1009 ();
 sg13g2_decap_8 FILLER_0_1016 ();
 sg13g2_decap_4 FILLER_0_1023 ();
 sg13g2_fill_2 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_fill_2 FILLER_1_91 ();
 sg13g2_fill_1 FILLER_1_93 ();
 sg13g2_fill_2 FILLER_1_103 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_fill_2 FILLER_1_147 ();
 sg13g2_fill_1 FILLER_1_149 ();
 sg13g2_decap_8 FILLER_1_177 ();
 sg13g2_decap_8 FILLER_1_184 ();
 sg13g2_decap_8 FILLER_1_191 ();
 sg13g2_decap_8 FILLER_1_198 ();
 sg13g2_decap_4 FILLER_1_205 ();
 sg13g2_fill_1 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_fill_1 FILLER_1_238 ();
 sg13g2_fill_2 FILLER_1_295 ();
 sg13g2_fill_1 FILLER_1_297 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_decap_8 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_1_435 ();
 sg13g2_decap_8 FILLER_1_442 ();
 sg13g2_decap_8 FILLER_1_449 ();
 sg13g2_decap_8 FILLER_1_456 ();
 sg13g2_decap_8 FILLER_1_463 ();
 sg13g2_decap_8 FILLER_1_470 ();
 sg13g2_decap_8 FILLER_1_477 ();
 sg13g2_decap_8 FILLER_1_484 ();
 sg13g2_decap_8 FILLER_1_491 ();
 sg13g2_decap_8 FILLER_1_498 ();
 sg13g2_decap_8 FILLER_1_505 ();
 sg13g2_decap_8 FILLER_1_512 ();
 sg13g2_decap_8 FILLER_1_519 ();
 sg13g2_decap_8 FILLER_1_526 ();
 sg13g2_decap_8 FILLER_1_533 ();
 sg13g2_decap_8 FILLER_1_540 ();
 sg13g2_decap_8 FILLER_1_547 ();
 sg13g2_decap_8 FILLER_1_554 ();
 sg13g2_decap_8 FILLER_1_561 ();
 sg13g2_decap_8 FILLER_1_568 ();
 sg13g2_decap_8 FILLER_1_575 ();
 sg13g2_decap_8 FILLER_1_582 ();
 sg13g2_decap_8 FILLER_1_589 ();
 sg13g2_decap_8 FILLER_1_596 ();
 sg13g2_decap_8 FILLER_1_603 ();
 sg13g2_decap_8 FILLER_1_610 ();
 sg13g2_decap_8 FILLER_1_617 ();
 sg13g2_decap_8 FILLER_1_624 ();
 sg13g2_decap_8 FILLER_1_631 ();
 sg13g2_decap_8 FILLER_1_638 ();
 sg13g2_decap_8 FILLER_1_645 ();
 sg13g2_decap_8 FILLER_1_652 ();
 sg13g2_decap_8 FILLER_1_659 ();
 sg13g2_decap_8 FILLER_1_666 ();
 sg13g2_decap_8 FILLER_1_673 ();
 sg13g2_decap_8 FILLER_1_680 ();
 sg13g2_decap_8 FILLER_1_687 ();
 sg13g2_decap_8 FILLER_1_694 ();
 sg13g2_decap_8 FILLER_1_701 ();
 sg13g2_decap_8 FILLER_1_708 ();
 sg13g2_decap_8 FILLER_1_715 ();
 sg13g2_decap_8 FILLER_1_722 ();
 sg13g2_decap_8 FILLER_1_729 ();
 sg13g2_decap_8 FILLER_1_736 ();
 sg13g2_decap_8 FILLER_1_743 ();
 sg13g2_decap_8 FILLER_1_750 ();
 sg13g2_decap_8 FILLER_1_757 ();
 sg13g2_decap_8 FILLER_1_764 ();
 sg13g2_decap_8 FILLER_1_771 ();
 sg13g2_decap_8 FILLER_1_778 ();
 sg13g2_decap_8 FILLER_1_785 ();
 sg13g2_decap_8 FILLER_1_792 ();
 sg13g2_decap_8 FILLER_1_799 ();
 sg13g2_decap_8 FILLER_1_806 ();
 sg13g2_decap_8 FILLER_1_813 ();
 sg13g2_decap_8 FILLER_1_820 ();
 sg13g2_decap_8 FILLER_1_827 ();
 sg13g2_decap_8 FILLER_1_834 ();
 sg13g2_decap_8 FILLER_1_841 ();
 sg13g2_decap_8 FILLER_1_848 ();
 sg13g2_decap_8 FILLER_1_855 ();
 sg13g2_decap_8 FILLER_1_862 ();
 sg13g2_decap_8 FILLER_1_869 ();
 sg13g2_decap_8 FILLER_1_876 ();
 sg13g2_decap_8 FILLER_1_883 ();
 sg13g2_decap_8 FILLER_1_890 ();
 sg13g2_decap_8 FILLER_1_897 ();
 sg13g2_decap_8 FILLER_1_904 ();
 sg13g2_decap_8 FILLER_1_911 ();
 sg13g2_decap_8 FILLER_1_918 ();
 sg13g2_decap_8 FILLER_1_925 ();
 sg13g2_decap_8 FILLER_1_932 ();
 sg13g2_decap_8 FILLER_1_939 ();
 sg13g2_decap_8 FILLER_1_946 ();
 sg13g2_decap_8 FILLER_1_953 ();
 sg13g2_decap_8 FILLER_1_960 ();
 sg13g2_decap_8 FILLER_1_967 ();
 sg13g2_decap_8 FILLER_1_974 ();
 sg13g2_decap_8 FILLER_1_981 ();
 sg13g2_decap_8 FILLER_1_988 ();
 sg13g2_decap_8 FILLER_1_995 ();
 sg13g2_decap_8 FILLER_1_1002 ();
 sg13g2_decap_8 FILLER_1_1009 ();
 sg13g2_decap_8 FILLER_1_1016 ();
 sg13g2_decap_4 FILLER_1_1023 ();
 sg13g2_fill_2 FILLER_1_1027 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_fill_2 FILLER_2_53 ();
 sg13g2_fill_1 FILLER_2_55 ();
 sg13g2_decap_8 FILLER_2_69 ();
 sg13g2_fill_1 FILLER_2_76 ();
 sg13g2_fill_2 FILLER_2_85 ();
 sg13g2_fill_1 FILLER_2_87 ();
 sg13g2_decap_4 FILLER_2_121 ();
 sg13g2_fill_2 FILLER_2_125 ();
 sg13g2_fill_2 FILLER_2_154 ();
 sg13g2_fill_1 FILLER_2_156 ();
 sg13g2_fill_1 FILLER_2_172 ();
 sg13g2_decap_4 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_190 ();
 sg13g2_decap_4 FILLER_2_197 ();
 sg13g2_fill_2 FILLER_2_218 ();
 sg13g2_fill_1 FILLER_2_220 ();
 sg13g2_fill_1 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_decap_8 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_2_436 ();
 sg13g2_decap_8 FILLER_2_443 ();
 sg13g2_decap_8 FILLER_2_450 ();
 sg13g2_decap_8 FILLER_2_457 ();
 sg13g2_decap_8 FILLER_2_464 ();
 sg13g2_decap_8 FILLER_2_471 ();
 sg13g2_decap_8 FILLER_2_478 ();
 sg13g2_decap_8 FILLER_2_485 ();
 sg13g2_decap_8 FILLER_2_492 ();
 sg13g2_decap_8 FILLER_2_499 ();
 sg13g2_decap_8 FILLER_2_506 ();
 sg13g2_decap_8 FILLER_2_513 ();
 sg13g2_decap_8 FILLER_2_520 ();
 sg13g2_decap_8 FILLER_2_527 ();
 sg13g2_decap_8 FILLER_2_534 ();
 sg13g2_decap_8 FILLER_2_541 ();
 sg13g2_decap_8 FILLER_2_548 ();
 sg13g2_decap_8 FILLER_2_555 ();
 sg13g2_decap_8 FILLER_2_562 ();
 sg13g2_decap_8 FILLER_2_569 ();
 sg13g2_decap_8 FILLER_2_576 ();
 sg13g2_decap_8 FILLER_2_583 ();
 sg13g2_decap_8 FILLER_2_590 ();
 sg13g2_decap_8 FILLER_2_597 ();
 sg13g2_decap_8 FILLER_2_604 ();
 sg13g2_decap_8 FILLER_2_611 ();
 sg13g2_decap_8 FILLER_2_618 ();
 sg13g2_decap_8 FILLER_2_625 ();
 sg13g2_decap_8 FILLER_2_632 ();
 sg13g2_decap_8 FILLER_2_639 ();
 sg13g2_decap_8 FILLER_2_646 ();
 sg13g2_decap_8 FILLER_2_653 ();
 sg13g2_decap_8 FILLER_2_660 ();
 sg13g2_decap_8 FILLER_2_667 ();
 sg13g2_decap_8 FILLER_2_674 ();
 sg13g2_decap_8 FILLER_2_681 ();
 sg13g2_decap_8 FILLER_2_688 ();
 sg13g2_decap_8 FILLER_2_695 ();
 sg13g2_decap_8 FILLER_2_702 ();
 sg13g2_decap_8 FILLER_2_709 ();
 sg13g2_decap_8 FILLER_2_716 ();
 sg13g2_decap_8 FILLER_2_723 ();
 sg13g2_decap_8 FILLER_2_730 ();
 sg13g2_decap_8 FILLER_2_737 ();
 sg13g2_decap_8 FILLER_2_744 ();
 sg13g2_decap_8 FILLER_2_751 ();
 sg13g2_decap_8 FILLER_2_758 ();
 sg13g2_decap_8 FILLER_2_765 ();
 sg13g2_decap_8 FILLER_2_772 ();
 sg13g2_decap_8 FILLER_2_779 ();
 sg13g2_decap_8 FILLER_2_786 ();
 sg13g2_decap_8 FILLER_2_793 ();
 sg13g2_decap_8 FILLER_2_800 ();
 sg13g2_decap_8 FILLER_2_807 ();
 sg13g2_decap_8 FILLER_2_814 ();
 sg13g2_decap_8 FILLER_2_821 ();
 sg13g2_decap_8 FILLER_2_828 ();
 sg13g2_decap_8 FILLER_2_835 ();
 sg13g2_decap_8 FILLER_2_842 ();
 sg13g2_decap_8 FILLER_2_849 ();
 sg13g2_decap_8 FILLER_2_856 ();
 sg13g2_decap_8 FILLER_2_863 ();
 sg13g2_decap_8 FILLER_2_870 ();
 sg13g2_decap_8 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_2_884 ();
 sg13g2_decap_8 FILLER_2_891 ();
 sg13g2_decap_8 FILLER_2_898 ();
 sg13g2_decap_8 FILLER_2_905 ();
 sg13g2_decap_8 FILLER_2_912 ();
 sg13g2_decap_8 FILLER_2_919 ();
 sg13g2_decap_8 FILLER_2_926 ();
 sg13g2_decap_8 FILLER_2_933 ();
 sg13g2_decap_8 FILLER_2_940 ();
 sg13g2_decap_8 FILLER_2_947 ();
 sg13g2_decap_8 FILLER_2_954 ();
 sg13g2_decap_8 FILLER_2_961 ();
 sg13g2_decap_8 FILLER_2_968 ();
 sg13g2_decap_8 FILLER_2_975 ();
 sg13g2_decap_8 FILLER_2_982 ();
 sg13g2_decap_8 FILLER_2_989 ();
 sg13g2_decap_8 FILLER_2_996 ();
 sg13g2_decap_8 FILLER_2_1003 ();
 sg13g2_decap_8 FILLER_2_1010 ();
 sg13g2_decap_8 FILLER_2_1017 ();
 sg13g2_decap_4 FILLER_2_1024 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_4 FILLER_3_46 ();
 sg13g2_fill_2 FILLER_3_86 ();
 sg13g2_fill_1 FILLER_3_88 ();
 sg13g2_fill_2 FILLER_3_105 ();
 sg13g2_fill_1 FILLER_3_107 ();
 sg13g2_fill_2 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_136 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_160 ();
 sg13g2_fill_1 FILLER_3_167 ();
 sg13g2_decap_4 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_fill_2 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_decap_8 FILLER_3_334 ();
 sg13g2_decap_8 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_8 FILLER_3_404 ();
 sg13g2_decap_8 FILLER_3_411 ();
 sg13g2_decap_8 FILLER_3_418 ();
 sg13g2_decap_8 FILLER_3_425 ();
 sg13g2_decap_8 FILLER_3_432 ();
 sg13g2_decap_8 FILLER_3_439 ();
 sg13g2_decap_8 FILLER_3_446 ();
 sg13g2_decap_8 FILLER_3_453 ();
 sg13g2_decap_8 FILLER_3_460 ();
 sg13g2_decap_8 FILLER_3_467 ();
 sg13g2_decap_8 FILLER_3_474 ();
 sg13g2_decap_8 FILLER_3_481 ();
 sg13g2_decap_8 FILLER_3_488 ();
 sg13g2_decap_8 FILLER_3_495 ();
 sg13g2_decap_8 FILLER_3_502 ();
 sg13g2_decap_8 FILLER_3_509 ();
 sg13g2_decap_8 FILLER_3_516 ();
 sg13g2_decap_8 FILLER_3_523 ();
 sg13g2_decap_8 FILLER_3_530 ();
 sg13g2_decap_8 FILLER_3_537 ();
 sg13g2_decap_8 FILLER_3_544 ();
 sg13g2_decap_8 FILLER_3_551 ();
 sg13g2_decap_8 FILLER_3_558 ();
 sg13g2_decap_8 FILLER_3_565 ();
 sg13g2_decap_8 FILLER_3_572 ();
 sg13g2_decap_8 FILLER_3_579 ();
 sg13g2_decap_8 FILLER_3_586 ();
 sg13g2_decap_8 FILLER_3_593 ();
 sg13g2_decap_8 FILLER_3_600 ();
 sg13g2_decap_8 FILLER_3_607 ();
 sg13g2_decap_8 FILLER_3_614 ();
 sg13g2_decap_8 FILLER_3_621 ();
 sg13g2_decap_8 FILLER_3_628 ();
 sg13g2_decap_8 FILLER_3_635 ();
 sg13g2_decap_8 FILLER_3_642 ();
 sg13g2_decap_8 FILLER_3_649 ();
 sg13g2_decap_8 FILLER_3_656 ();
 sg13g2_decap_8 FILLER_3_663 ();
 sg13g2_decap_8 FILLER_3_670 ();
 sg13g2_decap_8 FILLER_3_677 ();
 sg13g2_decap_8 FILLER_3_684 ();
 sg13g2_decap_8 FILLER_3_691 ();
 sg13g2_decap_8 FILLER_3_698 ();
 sg13g2_decap_8 FILLER_3_705 ();
 sg13g2_decap_8 FILLER_3_712 ();
 sg13g2_decap_8 FILLER_3_719 ();
 sg13g2_decap_8 FILLER_3_726 ();
 sg13g2_decap_8 FILLER_3_733 ();
 sg13g2_decap_8 FILLER_3_740 ();
 sg13g2_decap_8 FILLER_3_747 ();
 sg13g2_decap_8 FILLER_3_754 ();
 sg13g2_decap_8 FILLER_3_761 ();
 sg13g2_decap_8 FILLER_3_768 ();
 sg13g2_decap_8 FILLER_3_775 ();
 sg13g2_decap_8 FILLER_3_782 ();
 sg13g2_decap_8 FILLER_3_789 ();
 sg13g2_decap_8 FILLER_3_796 ();
 sg13g2_decap_8 FILLER_3_803 ();
 sg13g2_decap_8 FILLER_3_810 ();
 sg13g2_decap_8 FILLER_3_817 ();
 sg13g2_decap_8 FILLER_3_824 ();
 sg13g2_decap_8 FILLER_3_831 ();
 sg13g2_decap_8 FILLER_3_838 ();
 sg13g2_decap_8 FILLER_3_845 ();
 sg13g2_decap_8 FILLER_3_852 ();
 sg13g2_decap_8 FILLER_3_859 ();
 sg13g2_decap_8 FILLER_3_866 ();
 sg13g2_decap_8 FILLER_3_873 ();
 sg13g2_decap_8 FILLER_3_880 ();
 sg13g2_decap_8 FILLER_3_887 ();
 sg13g2_decap_8 FILLER_3_894 ();
 sg13g2_decap_8 FILLER_3_901 ();
 sg13g2_decap_8 FILLER_3_908 ();
 sg13g2_decap_8 FILLER_3_915 ();
 sg13g2_decap_8 FILLER_3_922 ();
 sg13g2_decap_8 FILLER_3_929 ();
 sg13g2_decap_8 FILLER_3_936 ();
 sg13g2_decap_8 FILLER_3_943 ();
 sg13g2_decap_8 FILLER_3_950 ();
 sg13g2_decap_8 FILLER_3_957 ();
 sg13g2_decap_8 FILLER_3_964 ();
 sg13g2_decap_8 FILLER_3_971 ();
 sg13g2_decap_8 FILLER_3_978 ();
 sg13g2_decap_8 FILLER_3_985 ();
 sg13g2_decap_8 FILLER_3_992 ();
 sg13g2_decap_8 FILLER_3_999 ();
 sg13g2_decap_8 FILLER_3_1006 ();
 sg13g2_decap_8 FILLER_3_1013 ();
 sg13g2_decap_8 FILLER_3_1020 ();
 sg13g2_fill_2 FILLER_3_1027 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_fill_2 FILLER_4_25 ();
 sg13g2_fill_1 FILLER_4_27 ();
 sg13g2_fill_2 FILLER_4_56 ();
 sg13g2_decap_4 FILLER_4_96 ();
 sg13g2_fill_2 FILLER_4_100 ();
 sg13g2_decap_8 FILLER_4_244 ();
 sg13g2_decap_4 FILLER_4_251 ();
 sg13g2_fill_2 FILLER_4_277 ();
 sg13g2_fill_1 FILLER_4_279 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_349 ();
 sg13g2_decap_8 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_8 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_4_412 ();
 sg13g2_decap_8 FILLER_4_419 ();
 sg13g2_decap_8 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_4_433 ();
 sg13g2_decap_8 FILLER_4_440 ();
 sg13g2_decap_8 FILLER_4_447 ();
 sg13g2_decap_8 FILLER_4_454 ();
 sg13g2_decap_8 FILLER_4_461 ();
 sg13g2_decap_8 FILLER_4_468 ();
 sg13g2_decap_8 FILLER_4_475 ();
 sg13g2_decap_8 FILLER_4_482 ();
 sg13g2_decap_8 FILLER_4_489 ();
 sg13g2_decap_8 FILLER_4_496 ();
 sg13g2_decap_8 FILLER_4_503 ();
 sg13g2_decap_8 FILLER_4_510 ();
 sg13g2_decap_8 FILLER_4_517 ();
 sg13g2_decap_8 FILLER_4_524 ();
 sg13g2_decap_8 FILLER_4_531 ();
 sg13g2_decap_8 FILLER_4_538 ();
 sg13g2_decap_8 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_552 ();
 sg13g2_decap_8 FILLER_4_559 ();
 sg13g2_decap_8 FILLER_4_566 ();
 sg13g2_decap_8 FILLER_4_573 ();
 sg13g2_decap_8 FILLER_4_580 ();
 sg13g2_decap_8 FILLER_4_587 ();
 sg13g2_decap_8 FILLER_4_594 ();
 sg13g2_decap_8 FILLER_4_601 ();
 sg13g2_decap_8 FILLER_4_608 ();
 sg13g2_decap_8 FILLER_4_615 ();
 sg13g2_decap_8 FILLER_4_622 ();
 sg13g2_decap_8 FILLER_4_629 ();
 sg13g2_decap_8 FILLER_4_636 ();
 sg13g2_decap_8 FILLER_4_643 ();
 sg13g2_decap_8 FILLER_4_650 ();
 sg13g2_decap_8 FILLER_4_657 ();
 sg13g2_decap_8 FILLER_4_664 ();
 sg13g2_decap_8 FILLER_4_671 ();
 sg13g2_decap_8 FILLER_4_678 ();
 sg13g2_decap_8 FILLER_4_685 ();
 sg13g2_decap_8 FILLER_4_692 ();
 sg13g2_decap_8 FILLER_4_699 ();
 sg13g2_decap_8 FILLER_4_706 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_decap_8 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_734 ();
 sg13g2_decap_8 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_748 ();
 sg13g2_decap_8 FILLER_4_755 ();
 sg13g2_decap_8 FILLER_4_762 ();
 sg13g2_decap_8 FILLER_4_769 ();
 sg13g2_decap_8 FILLER_4_776 ();
 sg13g2_decap_8 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_797 ();
 sg13g2_decap_8 FILLER_4_804 ();
 sg13g2_decap_8 FILLER_4_811 ();
 sg13g2_decap_8 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_825 ();
 sg13g2_decap_8 FILLER_4_832 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_853 ();
 sg13g2_decap_8 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_874 ();
 sg13g2_decap_8 FILLER_4_881 ();
 sg13g2_decap_8 FILLER_4_888 ();
 sg13g2_decap_8 FILLER_4_895 ();
 sg13g2_decap_8 FILLER_4_902 ();
 sg13g2_decap_8 FILLER_4_909 ();
 sg13g2_decap_8 FILLER_4_916 ();
 sg13g2_decap_8 FILLER_4_923 ();
 sg13g2_decap_8 FILLER_4_930 ();
 sg13g2_decap_8 FILLER_4_937 ();
 sg13g2_decap_8 FILLER_4_944 ();
 sg13g2_decap_8 FILLER_4_951 ();
 sg13g2_decap_8 FILLER_4_958 ();
 sg13g2_decap_8 FILLER_4_965 ();
 sg13g2_decap_8 FILLER_4_972 ();
 sg13g2_decap_8 FILLER_4_979 ();
 sg13g2_decap_8 FILLER_4_986 ();
 sg13g2_decap_8 FILLER_4_993 ();
 sg13g2_decap_8 FILLER_4_1000 ();
 sg13g2_decap_8 FILLER_4_1007 ();
 sg13g2_decap_8 FILLER_4_1014 ();
 sg13g2_decap_8 FILLER_4_1021 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_fill_1 FILLER_5_32 ();
 sg13g2_fill_2 FILLER_5_51 ();
 sg13g2_fill_2 FILLER_5_112 ();
 sg13g2_fill_1 FILLER_5_114 ();
 sg13g2_fill_1 FILLER_5_135 ();
 sg13g2_fill_1 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_1 FILLER_5_263 ();
 sg13g2_fill_1 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_5_430 ();
 sg13g2_decap_8 FILLER_5_437 ();
 sg13g2_decap_8 FILLER_5_444 ();
 sg13g2_decap_8 FILLER_5_451 ();
 sg13g2_decap_8 FILLER_5_458 ();
 sg13g2_decap_8 FILLER_5_465 ();
 sg13g2_decap_8 FILLER_5_472 ();
 sg13g2_decap_8 FILLER_5_479 ();
 sg13g2_decap_8 FILLER_5_486 ();
 sg13g2_decap_8 FILLER_5_493 ();
 sg13g2_decap_8 FILLER_5_500 ();
 sg13g2_decap_8 FILLER_5_507 ();
 sg13g2_decap_8 FILLER_5_514 ();
 sg13g2_decap_8 FILLER_5_521 ();
 sg13g2_decap_8 FILLER_5_528 ();
 sg13g2_decap_8 FILLER_5_535 ();
 sg13g2_decap_8 FILLER_5_542 ();
 sg13g2_decap_8 FILLER_5_549 ();
 sg13g2_decap_8 FILLER_5_556 ();
 sg13g2_decap_8 FILLER_5_563 ();
 sg13g2_decap_8 FILLER_5_570 ();
 sg13g2_decap_8 FILLER_5_577 ();
 sg13g2_decap_8 FILLER_5_584 ();
 sg13g2_decap_8 FILLER_5_591 ();
 sg13g2_decap_8 FILLER_5_598 ();
 sg13g2_decap_8 FILLER_5_605 ();
 sg13g2_decap_8 FILLER_5_612 ();
 sg13g2_decap_8 FILLER_5_619 ();
 sg13g2_decap_8 FILLER_5_626 ();
 sg13g2_decap_8 FILLER_5_633 ();
 sg13g2_decap_8 FILLER_5_640 ();
 sg13g2_decap_8 FILLER_5_647 ();
 sg13g2_decap_8 FILLER_5_654 ();
 sg13g2_decap_8 FILLER_5_661 ();
 sg13g2_decap_8 FILLER_5_668 ();
 sg13g2_decap_8 FILLER_5_675 ();
 sg13g2_decap_8 FILLER_5_682 ();
 sg13g2_decap_8 FILLER_5_689 ();
 sg13g2_decap_8 FILLER_5_696 ();
 sg13g2_decap_8 FILLER_5_703 ();
 sg13g2_decap_8 FILLER_5_710 ();
 sg13g2_decap_8 FILLER_5_717 ();
 sg13g2_decap_8 FILLER_5_724 ();
 sg13g2_decap_8 FILLER_5_731 ();
 sg13g2_decap_8 FILLER_5_738 ();
 sg13g2_decap_8 FILLER_5_745 ();
 sg13g2_decap_8 FILLER_5_752 ();
 sg13g2_decap_8 FILLER_5_759 ();
 sg13g2_decap_8 FILLER_5_766 ();
 sg13g2_decap_8 FILLER_5_773 ();
 sg13g2_decap_8 FILLER_5_780 ();
 sg13g2_decap_8 FILLER_5_787 ();
 sg13g2_decap_8 FILLER_5_794 ();
 sg13g2_decap_8 FILLER_5_801 ();
 sg13g2_decap_8 FILLER_5_808 ();
 sg13g2_decap_8 FILLER_5_815 ();
 sg13g2_decap_8 FILLER_5_822 ();
 sg13g2_decap_8 FILLER_5_829 ();
 sg13g2_decap_8 FILLER_5_836 ();
 sg13g2_decap_8 FILLER_5_843 ();
 sg13g2_decap_8 FILLER_5_850 ();
 sg13g2_decap_8 FILLER_5_857 ();
 sg13g2_decap_8 FILLER_5_864 ();
 sg13g2_decap_8 FILLER_5_871 ();
 sg13g2_decap_8 FILLER_5_878 ();
 sg13g2_decap_8 FILLER_5_885 ();
 sg13g2_decap_8 FILLER_5_892 ();
 sg13g2_decap_8 FILLER_5_899 ();
 sg13g2_decap_8 FILLER_5_906 ();
 sg13g2_decap_8 FILLER_5_913 ();
 sg13g2_decap_8 FILLER_5_920 ();
 sg13g2_decap_8 FILLER_5_927 ();
 sg13g2_decap_8 FILLER_5_934 ();
 sg13g2_decap_8 FILLER_5_941 ();
 sg13g2_decap_8 FILLER_5_948 ();
 sg13g2_decap_8 FILLER_5_955 ();
 sg13g2_decap_8 FILLER_5_962 ();
 sg13g2_decap_8 FILLER_5_969 ();
 sg13g2_decap_8 FILLER_5_976 ();
 sg13g2_decap_8 FILLER_5_983 ();
 sg13g2_decap_8 FILLER_5_990 ();
 sg13g2_decap_8 FILLER_5_997 ();
 sg13g2_decap_8 FILLER_5_1004 ();
 sg13g2_decap_8 FILLER_5_1011 ();
 sg13g2_decap_8 FILLER_5_1018 ();
 sg13g2_decap_4 FILLER_5_1025 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_fill_2 FILLER_6_32 ();
 sg13g2_fill_1 FILLER_6_34 ();
 sg13g2_fill_1 FILLER_6_56 ();
 sg13g2_fill_1 FILLER_6_93 ();
 sg13g2_fill_1 FILLER_6_108 ();
 sg13g2_fill_1 FILLER_6_119 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_fill_2 FILLER_6_172 ();
 sg13g2_fill_1 FILLER_6_174 ();
 sg13g2_fill_1 FILLER_6_179 ();
 sg13g2_fill_2 FILLER_6_208 ();
 sg13g2_fill_1 FILLER_6_210 ();
 sg13g2_fill_1 FILLER_6_239 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_decap_4 FILLER_6_269 ();
 sg13g2_decap_4 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_fill_2 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_8 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_6_412 ();
 sg13g2_decap_8 FILLER_6_419 ();
 sg13g2_decap_8 FILLER_6_426 ();
 sg13g2_decap_8 FILLER_6_433 ();
 sg13g2_decap_8 FILLER_6_440 ();
 sg13g2_decap_8 FILLER_6_447 ();
 sg13g2_decap_8 FILLER_6_454 ();
 sg13g2_decap_8 FILLER_6_461 ();
 sg13g2_decap_8 FILLER_6_468 ();
 sg13g2_decap_8 FILLER_6_475 ();
 sg13g2_decap_8 FILLER_6_482 ();
 sg13g2_decap_8 FILLER_6_489 ();
 sg13g2_decap_8 FILLER_6_496 ();
 sg13g2_decap_8 FILLER_6_503 ();
 sg13g2_decap_8 FILLER_6_510 ();
 sg13g2_decap_8 FILLER_6_517 ();
 sg13g2_decap_8 FILLER_6_524 ();
 sg13g2_decap_8 FILLER_6_531 ();
 sg13g2_decap_8 FILLER_6_538 ();
 sg13g2_decap_8 FILLER_6_545 ();
 sg13g2_decap_8 FILLER_6_552 ();
 sg13g2_decap_8 FILLER_6_559 ();
 sg13g2_decap_8 FILLER_6_566 ();
 sg13g2_decap_8 FILLER_6_573 ();
 sg13g2_decap_8 FILLER_6_580 ();
 sg13g2_decap_8 FILLER_6_587 ();
 sg13g2_decap_8 FILLER_6_594 ();
 sg13g2_decap_8 FILLER_6_601 ();
 sg13g2_decap_8 FILLER_6_608 ();
 sg13g2_decap_8 FILLER_6_615 ();
 sg13g2_decap_8 FILLER_6_622 ();
 sg13g2_decap_8 FILLER_6_629 ();
 sg13g2_decap_8 FILLER_6_636 ();
 sg13g2_decap_8 FILLER_6_643 ();
 sg13g2_decap_8 FILLER_6_650 ();
 sg13g2_decap_8 FILLER_6_657 ();
 sg13g2_decap_8 FILLER_6_664 ();
 sg13g2_decap_8 FILLER_6_671 ();
 sg13g2_decap_8 FILLER_6_678 ();
 sg13g2_decap_8 FILLER_6_685 ();
 sg13g2_decap_8 FILLER_6_692 ();
 sg13g2_decap_8 FILLER_6_699 ();
 sg13g2_decap_8 FILLER_6_706 ();
 sg13g2_decap_8 FILLER_6_713 ();
 sg13g2_decap_8 FILLER_6_720 ();
 sg13g2_decap_8 FILLER_6_727 ();
 sg13g2_decap_8 FILLER_6_734 ();
 sg13g2_decap_8 FILLER_6_741 ();
 sg13g2_decap_8 FILLER_6_748 ();
 sg13g2_decap_8 FILLER_6_755 ();
 sg13g2_decap_8 FILLER_6_762 ();
 sg13g2_decap_8 FILLER_6_769 ();
 sg13g2_decap_8 FILLER_6_776 ();
 sg13g2_decap_8 FILLER_6_783 ();
 sg13g2_decap_8 FILLER_6_790 ();
 sg13g2_decap_8 FILLER_6_797 ();
 sg13g2_decap_8 FILLER_6_804 ();
 sg13g2_decap_8 FILLER_6_811 ();
 sg13g2_decap_8 FILLER_6_818 ();
 sg13g2_decap_8 FILLER_6_825 ();
 sg13g2_decap_8 FILLER_6_832 ();
 sg13g2_decap_8 FILLER_6_839 ();
 sg13g2_decap_8 FILLER_6_846 ();
 sg13g2_decap_8 FILLER_6_853 ();
 sg13g2_decap_8 FILLER_6_860 ();
 sg13g2_decap_8 FILLER_6_867 ();
 sg13g2_decap_8 FILLER_6_874 ();
 sg13g2_decap_8 FILLER_6_881 ();
 sg13g2_decap_8 FILLER_6_888 ();
 sg13g2_decap_8 FILLER_6_895 ();
 sg13g2_decap_8 FILLER_6_902 ();
 sg13g2_decap_8 FILLER_6_909 ();
 sg13g2_decap_8 FILLER_6_916 ();
 sg13g2_decap_8 FILLER_6_923 ();
 sg13g2_decap_8 FILLER_6_930 ();
 sg13g2_decap_8 FILLER_6_937 ();
 sg13g2_decap_8 FILLER_6_944 ();
 sg13g2_decap_8 FILLER_6_951 ();
 sg13g2_decap_8 FILLER_6_958 ();
 sg13g2_decap_8 FILLER_6_965 ();
 sg13g2_decap_8 FILLER_6_972 ();
 sg13g2_decap_8 FILLER_6_979 ();
 sg13g2_decap_8 FILLER_6_986 ();
 sg13g2_decap_8 FILLER_6_993 ();
 sg13g2_decap_8 FILLER_6_1000 ();
 sg13g2_decap_8 FILLER_6_1007 ();
 sg13g2_decap_8 FILLER_6_1014 ();
 sg13g2_decap_8 FILLER_6_1021 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_4 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_77 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_121 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_135 ();
 sg13g2_fill_1 FILLER_7_144 ();
 sg13g2_fill_1 FILLER_7_184 ();
 sg13g2_fill_2 FILLER_7_193 ();
 sg13g2_fill_1 FILLER_7_195 ();
 sg13g2_fill_2 FILLER_7_209 ();
 sg13g2_decap_8 FILLER_7_278 ();
 sg13g2_fill_2 FILLER_7_285 ();
 sg13g2_fill_1 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_8 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_7_412 ();
 sg13g2_decap_8 FILLER_7_419 ();
 sg13g2_decap_8 FILLER_7_426 ();
 sg13g2_decap_8 FILLER_7_433 ();
 sg13g2_decap_8 FILLER_7_440 ();
 sg13g2_decap_8 FILLER_7_447 ();
 sg13g2_decap_8 FILLER_7_454 ();
 sg13g2_decap_8 FILLER_7_461 ();
 sg13g2_decap_8 FILLER_7_468 ();
 sg13g2_decap_8 FILLER_7_475 ();
 sg13g2_decap_8 FILLER_7_482 ();
 sg13g2_decap_8 FILLER_7_489 ();
 sg13g2_decap_8 FILLER_7_496 ();
 sg13g2_decap_8 FILLER_7_503 ();
 sg13g2_decap_8 FILLER_7_510 ();
 sg13g2_decap_8 FILLER_7_517 ();
 sg13g2_decap_8 FILLER_7_524 ();
 sg13g2_decap_8 FILLER_7_531 ();
 sg13g2_decap_8 FILLER_7_538 ();
 sg13g2_decap_8 FILLER_7_545 ();
 sg13g2_decap_8 FILLER_7_552 ();
 sg13g2_decap_8 FILLER_7_559 ();
 sg13g2_decap_8 FILLER_7_566 ();
 sg13g2_decap_8 FILLER_7_573 ();
 sg13g2_decap_8 FILLER_7_580 ();
 sg13g2_decap_8 FILLER_7_587 ();
 sg13g2_decap_8 FILLER_7_594 ();
 sg13g2_decap_8 FILLER_7_601 ();
 sg13g2_decap_8 FILLER_7_608 ();
 sg13g2_decap_8 FILLER_7_615 ();
 sg13g2_decap_8 FILLER_7_622 ();
 sg13g2_decap_8 FILLER_7_629 ();
 sg13g2_decap_8 FILLER_7_636 ();
 sg13g2_decap_8 FILLER_7_643 ();
 sg13g2_decap_8 FILLER_7_650 ();
 sg13g2_decap_8 FILLER_7_657 ();
 sg13g2_decap_8 FILLER_7_664 ();
 sg13g2_decap_8 FILLER_7_671 ();
 sg13g2_decap_8 FILLER_7_678 ();
 sg13g2_decap_8 FILLER_7_685 ();
 sg13g2_decap_8 FILLER_7_692 ();
 sg13g2_decap_8 FILLER_7_699 ();
 sg13g2_decap_8 FILLER_7_706 ();
 sg13g2_decap_8 FILLER_7_713 ();
 sg13g2_decap_8 FILLER_7_720 ();
 sg13g2_decap_8 FILLER_7_727 ();
 sg13g2_decap_8 FILLER_7_734 ();
 sg13g2_decap_8 FILLER_7_741 ();
 sg13g2_decap_8 FILLER_7_748 ();
 sg13g2_decap_8 FILLER_7_755 ();
 sg13g2_decap_8 FILLER_7_762 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_8 FILLER_7_804 ();
 sg13g2_decap_8 FILLER_7_811 ();
 sg13g2_decap_8 FILLER_7_818 ();
 sg13g2_decap_8 FILLER_7_825 ();
 sg13g2_decap_8 FILLER_7_832 ();
 sg13g2_decap_8 FILLER_7_839 ();
 sg13g2_decap_8 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_853 ();
 sg13g2_decap_8 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_7_867 ();
 sg13g2_decap_8 FILLER_7_874 ();
 sg13g2_decap_8 FILLER_7_881 ();
 sg13g2_decap_8 FILLER_7_888 ();
 sg13g2_decap_8 FILLER_7_895 ();
 sg13g2_decap_8 FILLER_7_902 ();
 sg13g2_decap_8 FILLER_7_909 ();
 sg13g2_decap_8 FILLER_7_916 ();
 sg13g2_decap_8 FILLER_7_923 ();
 sg13g2_decap_8 FILLER_7_930 ();
 sg13g2_decap_8 FILLER_7_937 ();
 sg13g2_decap_8 FILLER_7_944 ();
 sg13g2_decap_8 FILLER_7_951 ();
 sg13g2_decap_8 FILLER_7_958 ();
 sg13g2_decap_8 FILLER_7_965 ();
 sg13g2_decap_8 FILLER_7_972 ();
 sg13g2_decap_8 FILLER_7_979 ();
 sg13g2_decap_8 FILLER_7_986 ();
 sg13g2_decap_8 FILLER_7_993 ();
 sg13g2_decap_8 FILLER_7_1000 ();
 sg13g2_decap_8 FILLER_7_1007 ();
 sg13g2_decap_8 FILLER_7_1014 ();
 sg13g2_decap_8 FILLER_7_1021 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_fill_1 FILLER_8_46 ();
 sg13g2_fill_1 FILLER_8_74 ();
 sg13g2_fill_2 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_139 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_fill_2 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_190 ();
 sg13g2_fill_1 FILLER_8_231 ();
 sg13g2_fill_2 FILLER_8_253 ();
 sg13g2_fill_1 FILLER_8_255 ();
 sg13g2_decap_4 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_283 ();
 sg13g2_decap_8 FILLER_8_310 ();
 sg13g2_fill_1 FILLER_8_317 ();
 sg13g2_fill_1 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_334 ();
 sg13g2_fill_2 FILLER_8_341 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_fill_2 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_decap_8 FILLER_8_875 ();
 sg13g2_decap_8 FILLER_8_882 ();
 sg13g2_decap_8 FILLER_8_889 ();
 sg13g2_decap_8 FILLER_8_896 ();
 sg13g2_decap_8 FILLER_8_903 ();
 sg13g2_decap_8 FILLER_8_910 ();
 sg13g2_decap_8 FILLER_8_917 ();
 sg13g2_decap_8 FILLER_8_924 ();
 sg13g2_decap_8 FILLER_8_931 ();
 sg13g2_decap_8 FILLER_8_938 ();
 sg13g2_decap_8 FILLER_8_945 ();
 sg13g2_decap_8 FILLER_8_952 ();
 sg13g2_decap_8 FILLER_8_959 ();
 sg13g2_decap_8 FILLER_8_966 ();
 sg13g2_decap_8 FILLER_8_973 ();
 sg13g2_decap_8 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_987 ();
 sg13g2_decap_8 FILLER_8_994 ();
 sg13g2_decap_8 FILLER_8_1001 ();
 sg13g2_decap_8 FILLER_8_1008 ();
 sg13g2_decap_8 FILLER_8_1015 ();
 sg13g2_decap_8 FILLER_8_1022 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_4 FILLER_9_18 ();
 sg13g2_fill_1 FILLER_9_22 ();
 sg13g2_decap_4 FILLER_9_27 ();
 sg13g2_fill_2 FILLER_9_31 ();
 sg13g2_decap_4 FILLER_9_66 ();
 sg13g2_fill_1 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_fill_2 FILLER_9_109 ();
 sg13g2_fill_1 FILLER_9_111 ();
 sg13g2_fill_2 FILLER_9_132 ();
 sg13g2_fill_1 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_240 ();
 sg13g2_decap_4 FILLER_9_246 ();
 sg13g2_fill_1 FILLER_9_250 ();
 sg13g2_decap_4 FILLER_9_264 ();
 sg13g2_decap_4 FILLER_9_281 ();
 sg13g2_fill_1 FILLER_9_285 ();
 sg13g2_fill_1 FILLER_9_302 ();
 sg13g2_fill_1 FILLER_9_316 ();
 sg13g2_fill_1 FILLER_9_323 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_9_409 ();
 sg13g2_decap_8 FILLER_9_416 ();
 sg13g2_decap_8 FILLER_9_423 ();
 sg13g2_decap_8 FILLER_9_430 ();
 sg13g2_decap_8 FILLER_9_437 ();
 sg13g2_decap_8 FILLER_9_444 ();
 sg13g2_decap_8 FILLER_9_451 ();
 sg13g2_decap_8 FILLER_9_458 ();
 sg13g2_decap_8 FILLER_9_465 ();
 sg13g2_decap_8 FILLER_9_472 ();
 sg13g2_decap_8 FILLER_9_479 ();
 sg13g2_decap_8 FILLER_9_486 ();
 sg13g2_decap_8 FILLER_9_493 ();
 sg13g2_decap_8 FILLER_9_500 ();
 sg13g2_decap_8 FILLER_9_507 ();
 sg13g2_decap_8 FILLER_9_514 ();
 sg13g2_decap_8 FILLER_9_521 ();
 sg13g2_decap_8 FILLER_9_528 ();
 sg13g2_decap_8 FILLER_9_535 ();
 sg13g2_decap_8 FILLER_9_542 ();
 sg13g2_decap_8 FILLER_9_549 ();
 sg13g2_decap_8 FILLER_9_556 ();
 sg13g2_decap_8 FILLER_9_563 ();
 sg13g2_decap_8 FILLER_9_570 ();
 sg13g2_decap_8 FILLER_9_577 ();
 sg13g2_decap_8 FILLER_9_584 ();
 sg13g2_decap_8 FILLER_9_591 ();
 sg13g2_decap_8 FILLER_9_598 ();
 sg13g2_decap_8 FILLER_9_605 ();
 sg13g2_decap_8 FILLER_9_612 ();
 sg13g2_decap_8 FILLER_9_619 ();
 sg13g2_decap_8 FILLER_9_626 ();
 sg13g2_decap_8 FILLER_9_633 ();
 sg13g2_decap_8 FILLER_9_640 ();
 sg13g2_decap_8 FILLER_9_647 ();
 sg13g2_decap_8 FILLER_9_654 ();
 sg13g2_decap_8 FILLER_9_661 ();
 sg13g2_decap_8 FILLER_9_668 ();
 sg13g2_decap_8 FILLER_9_675 ();
 sg13g2_decap_8 FILLER_9_682 ();
 sg13g2_decap_8 FILLER_9_689 ();
 sg13g2_decap_8 FILLER_9_696 ();
 sg13g2_decap_8 FILLER_9_703 ();
 sg13g2_decap_8 FILLER_9_710 ();
 sg13g2_decap_8 FILLER_9_717 ();
 sg13g2_decap_8 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_731 ();
 sg13g2_decap_8 FILLER_9_738 ();
 sg13g2_decap_8 FILLER_9_745 ();
 sg13g2_decap_8 FILLER_9_752 ();
 sg13g2_decap_8 FILLER_9_759 ();
 sg13g2_decap_8 FILLER_9_766 ();
 sg13g2_decap_8 FILLER_9_773 ();
 sg13g2_decap_8 FILLER_9_780 ();
 sg13g2_decap_8 FILLER_9_787 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_decap_8 FILLER_9_801 ();
 sg13g2_decap_8 FILLER_9_808 ();
 sg13g2_decap_8 FILLER_9_815 ();
 sg13g2_decap_8 FILLER_9_822 ();
 sg13g2_decap_8 FILLER_9_829 ();
 sg13g2_decap_8 FILLER_9_836 ();
 sg13g2_decap_8 FILLER_9_843 ();
 sg13g2_decap_8 FILLER_9_850 ();
 sg13g2_decap_8 FILLER_9_857 ();
 sg13g2_decap_8 FILLER_9_864 ();
 sg13g2_decap_8 FILLER_9_871 ();
 sg13g2_decap_8 FILLER_9_878 ();
 sg13g2_decap_8 FILLER_9_885 ();
 sg13g2_decap_8 FILLER_9_892 ();
 sg13g2_decap_8 FILLER_9_899 ();
 sg13g2_decap_8 FILLER_9_906 ();
 sg13g2_decap_8 FILLER_9_913 ();
 sg13g2_decap_8 FILLER_9_920 ();
 sg13g2_decap_8 FILLER_9_927 ();
 sg13g2_decap_8 FILLER_9_934 ();
 sg13g2_decap_8 FILLER_9_941 ();
 sg13g2_decap_8 FILLER_9_948 ();
 sg13g2_decap_8 FILLER_9_955 ();
 sg13g2_decap_8 FILLER_9_962 ();
 sg13g2_decap_8 FILLER_9_969 ();
 sg13g2_decap_8 FILLER_9_976 ();
 sg13g2_decap_8 FILLER_9_983 ();
 sg13g2_decap_8 FILLER_9_990 ();
 sg13g2_decap_8 FILLER_9_997 ();
 sg13g2_decap_8 FILLER_9_1004 ();
 sg13g2_decap_8 FILLER_9_1011 ();
 sg13g2_decap_8 FILLER_9_1018 ();
 sg13g2_decap_4 FILLER_9_1025 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_4 FILLER_10_25 ();
 sg13g2_fill_2 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_90 ();
 sg13g2_fill_2 FILLER_10_106 ();
 sg13g2_fill_2 FILLER_10_144 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_185 ();
 sg13g2_decap_8 FILLER_10_192 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_decap_4 FILLER_10_228 ();
 sg13g2_fill_2 FILLER_10_247 ();
 sg13g2_fill_1 FILLER_10_249 ();
 sg13g2_fill_1 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_4 FILLER_10_287 ();
 sg13g2_fill_2 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_316 ();
 sg13g2_fill_1 FILLER_10_341 ();
 sg13g2_fill_2 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_424 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_8 FILLER_10_438 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_decap_8 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_decap_8 FILLER_10_466 ();
 sg13g2_decap_8 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_decap_8 FILLER_10_501 ();
 sg13g2_decap_8 FILLER_10_508 ();
 sg13g2_decap_8 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_522 ();
 sg13g2_decap_8 FILLER_10_529 ();
 sg13g2_decap_8 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_550 ();
 sg13g2_decap_8 FILLER_10_557 ();
 sg13g2_decap_8 FILLER_10_564 ();
 sg13g2_decap_8 FILLER_10_571 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_decap_8 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_669 ();
 sg13g2_decap_8 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_683 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_872 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_decap_8 FILLER_10_886 ();
 sg13g2_decap_8 FILLER_10_893 ();
 sg13g2_decap_8 FILLER_10_900 ();
 sg13g2_decap_8 FILLER_10_907 ();
 sg13g2_decap_8 FILLER_10_914 ();
 sg13g2_decap_8 FILLER_10_921 ();
 sg13g2_decap_8 FILLER_10_928 ();
 sg13g2_decap_8 FILLER_10_935 ();
 sg13g2_decap_8 FILLER_10_942 ();
 sg13g2_decap_8 FILLER_10_949 ();
 sg13g2_decap_8 FILLER_10_956 ();
 sg13g2_decap_8 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_970 ();
 sg13g2_decap_8 FILLER_10_977 ();
 sg13g2_decap_8 FILLER_10_984 ();
 sg13g2_decap_8 FILLER_10_991 ();
 sg13g2_decap_8 FILLER_10_998 ();
 sg13g2_decap_8 FILLER_10_1005 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_fill_2 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_fill_2 FILLER_11_32 ();
 sg13g2_decap_8 FILLER_11_38 ();
 sg13g2_decap_4 FILLER_11_45 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_95 ();
 sg13g2_decap_4 FILLER_11_104 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_169 ();
 sg13g2_decap_8 FILLER_11_192 ();
 sg13g2_decap_4 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_203 ();
 sg13g2_decap_4 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_226 ();
 sg13g2_fill_1 FILLER_11_243 ();
 sg13g2_fill_2 FILLER_11_254 ();
 sg13g2_decap_8 FILLER_11_260 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_fill_2 FILLER_11_274 ();
 sg13g2_fill_1 FILLER_11_276 ();
 sg13g2_fill_1 FILLER_11_286 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_fill_2 FILLER_11_322 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_330 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_fill_2 FILLER_11_369 ();
 sg13g2_fill_2 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_decap_8 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_11_435 ();
 sg13g2_decap_8 FILLER_11_442 ();
 sg13g2_decap_8 FILLER_11_449 ();
 sg13g2_decap_8 FILLER_11_456 ();
 sg13g2_decap_8 FILLER_11_463 ();
 sg13g2_decap_8 FILLER_11_470 ();
 sg13g2_decap_8 FILLER_11_477 ();
 sg13g2_decap_8 FILLER_11_484 ();
 sg13g2_decap_8 FILLER_11_491 ();
 sg13g2_decap_8 FILLER_11_498 ();
 sg13g2_decap_8 FILLER_11_505 ();
 sg13g2_decap_8 FILLER_11_512 ();
 sg13g2_decap_8 FILLER_11_519 ();
 sg13g2_decap_8 FILLER_11_526 ();
 sg13g2_decap_8 FILLER_11_533 ();
 sg13g2_decap_8 FILLER_11_540 ();
 sg13g2_decap_8 FILLER_11_547 ();
 sg13g2_decap_8 FILLER_11_554 ();
 sg13g2_decap_8 FILLER_11_561 ();
 sg13g2_decap_8 FILLER_11_568 ();
 sg13g2_decap_8 FILLER_11_575 ();
 sg13g2_decap_8 FILLER_11_582 ();
 sg13g2_decap_8 FILLER_11_589 ();
 sg13g2_decap_8 FILLER_11_596 ();
 sg13g2_decap_8 FILLER_11_603 ();
 sg13g2_decap_8 FILLER_11_610 ();
 sg13g2_decap_8 FILLER_11_617 ();
 sg13g2_decap_8 FILLER_11_624 ();
 sg13g2_decap_8 FILLER_11_631 ();
 sg13g2_decap_8 FILLER_11_638 ();
 sg13g2_decap_8 FILLER_11_645 ();
 sg13g2_decap_8 FILLER_11_652 ();
 sg13g2_decap_8 FILLER_11_659 ();
 sg13g2_decap_8 FILLER_11_666 ();
 sg13g2_decap_8 FILLER_11_673 ();
 sg13g2_decap_8 FILLER_11_680 ();
 sg13g2_decap_8 FILLER_11_687 ();
 sg13g2_decap_8 FILLER_11_694 ();
 sg13g2_decap_8 FILLER_11_701 ();
 sg13g2_decap_8 FILLER_11_708 ();
 sg13g2_decap_8 FILLER_11_715 ();
 sg13g2_decap_8 FILLER_11_722 ();
 sg13g2_decap_8 FILLER_11_729 ();
 sg13g2_decap_8 FILLER_11_736 ();
 sg13g2_decap_8 FILLER_11_743 ();
 sg13g2_decap_8 FILLER_11_750 ();
 sg13g2_decap_8 FILLER_11_757 ();
 sg13g2_decap_8 FILLER_11_764 ();
 sg13g2_decap_8 FILLER_11_771 ();
 sg13g2_decap_8 FILLER_11_778 ();
 sg13g2_decap_8 FILLER_11_785 ();
 sg13g2_decap_8 FILLER_11_792 ();
 sg13g2_decap_8 FILLER_11_799 ();
 sg13g2_decap_8 FILLER_11_806 ();
 sg13g2_decap_8 FILLER_11_813 ();
 sg13g2_decap_8 FILLER_11_820 ();
 sg13g2_decap_8 FILLER_11_827 ();
 sg13g2_decap_8 FILLER_11_834 ();
 sg13g2_decap_8 FILLER_11_841 ();
 sg13g2_decap_8 FILLER_11_848 ();
 sg13g2_decap_8 FILLER_11_855 ();
 sg13g2_decap_8 FILLER_11_862 ();
 sg13g2_decap_8 FILLER_11_869 ();
 sg13g2_decap_8 FILLER_11_876 ();
 sg13g2_decap_8 FILLER_11_883 ();
 sg13g2_decap_8 FILLER_11_890 ();
 sg13g2_decap_8 FILLER_11_897 ();
 sg13g2_decap_8 FILLER_11_904 ();
 sg13g2_decap_8 FILLER_11_911 ();
 sg13g2_decap_8 FILLER_11_918 ();
 sg13g2_decap_8 FILLER_11_925 ();
 sg13g2_decap_8 FILLER_11_932 ();
 sg13g2_decap_8 FILLER_11_939 ();
 sg13g2_decap_8 FILLER_11_946 ();
 sg13g2_decap_8 FILLER_11_953 ();
 sg13g2_decap_8 FILLER_11_960 ();
 sg13g2_decap_8 FILLER_11_967 ();
 sg13g2_decap_8 FILLER_11_974 ();
 sg13g2_decap_8 FILLER_11_981 ();
 sg13g2_decap_8 FILLER_11_988 ();
 sg13g2_decap_8 FILLER_11_995 ();
 sg13g2_decap_8 FILLER_11_1002 ();
 sg13g2_decap_8 FILLER_11_1009 ();
 sg13g2_decap_8 FILLER_11_1016 ();
 sg13g2_decap_4 FILLER_11_1023 ();
 sg13g2_fill_2 FILLER_11_1027 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_46 ();
 sg13g2_fill_2 FILLER_12_53 ();
 sg13g2_fill_1 FILLER_12_55 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_159 ();
 sg13g2_fill_2 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_279 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_fill_1 FILLER_12_293 ();
 sg13g2_fill_2 FILLER_12_312 ();
 sg13g2_decap_4 FILLER_12_322 ();
 sg13g2_fill_2 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_4 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_8 FILLER_12_425 ();
 sg13g2_decap_8 FILLER_12_432 ();
 sg13g2_decap_8 FILLER_12_439 ();
 sg13g2_decap_8 FILLER_12_446 ();
 sg13g2_decap_8 FILLER_12_453 ();
 sg13g2_decap_8 FILLER_12_460 ();
 sg13g2_decap_8 FILLER_12_467 ();
 sg13g2_decap_8 FILLER_12_474 ();
 sg13g2_decap_8 FILLER_12_481 ();
 sg13g2_decap_8 FILLER_12_488 ();
 sg13g2_decap_8 FILLER_12_495 ();
 sg13g2_decap_8 FILLER_12_502 ();
 sg13g2_decap_8 FILLER_12_509 ();
 sg13g2_decap_8 FILLER_12_516 ();
 sg13g2_decap_8 FILLER_12_523 ();
 sg13g2_decap_8 FILLER_12_530 ();
 sg13g2_decap_8 FILLER_12_537 ();
 sg13g2_decap_8 FILLER_12_544 ();
 sg13g2_decap_8 FILLER_12_551 ();
 sg13g2_decap_8 FILLER_12_558 ();
 sg13g2_decap_8 FILLER_12_565 ();
 sg13g2_decap_8 FILLER_12_572 ();
 sg13g2_decap_8 FILLER_12_579 ();
 sg13g2_decap_8 FILLER_12_586 ();
 sg13g2_decap_8 FILLER_12_593 ();
 sg13g2_decap_8 FILLER_12_600 ();
 sg13g2_decap_8 FILLER_12_607 ();
 sg13g2_decap_8 FILLER_12_614 ();
 sg13g2_decap_8 FILLER_12_621 ();
 sg13g2_decap_8 FILLER_12_628 ();
 sg13g2_decap_8 FILLER_12_635 ();
 sg13g2_decap_8 FILLER_12_642 ();
 sg13g2_decap_8 FILLER_12_649 ();
 sg13g2_decap_8 FILLER_12_656 ();
 sg13g2_decap_8 FILLER_12_663 ();
 sg13g2_decap_8 FILLER_12_670 ();
 sg13g2_decap_8 FILLER_12_677 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_decap_8 FILLER_12_691 ();
 sg13g2_decap_8 FILLER_12_698 ();
 sg13g2_decap_8 FILLER_12_705 ();
 sg13g2_decap_8 FILLER_12_712 ();
 sg13g2_decap_8 FILLER_12_719 ();
 sg13g2_decap_8 FILLER_12_726 ();
 sg13g2_decap_8 FILLER_12_733 ();
 sg13g2_decap_8 FILLER_12_740 ();
 sg13g2_decap_8 FILLER_12_747 ();
 sg13g2_decap_8 FILLER_12_754 ();
 sg13g2_decap_8 FILLER_12_761 ();
 sg13g2_decap_8 FILLER_12_768 ();
 sg13g2_decap_8 FILLER_12_775 ();
 sg13g2_decap_8 FILLER_12_782 ();
 sg13g2_decap_8 FILLER_12_789 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_decap_8 FILLER_12_803 ();
 sg13g2_decap_8 FILLER_12_810 ();
 sg13g2_decap_8 FILLER_12_817 ();
 sg13g2_decap_8 FILLER_12_824 ();
 sg13g2_decap_8 FILLER_12_831 ();
 sg13g2_decap_8 FILLER_12_838 ();
 sg13g2_decap_8 FILLER_12_845 ();
 sg13g2_decap_8 FILLER_12_852 ();
 sg13g2_decap_8 FILLER_12_859 ();
 sg13g2_decap_8 FILLER_12_866 ();
 sg13g2_decap_8 FILLER_12_873 ();
 sg13g2_decap_8 FILLER_12_880 ();
 sg13g2_decap_8 FILLER_12_887 ();
 sg13g2_decap_8 FILLER_12_894 ();
 sg13g2_decap_8 FILLER_12_901 ();
 sg13g2_decap_8 FILLER_12_908 ();
 sg13g2_decap_8 FILLER_12_915 ();
 sg13g2_decap_8 FILLER_12_922 ();
 sg13g2_decap_8 FILLER_12_929 ();
 sg13g2_decap_8 FILLER_12_936 ();
 sg13g2_decap_8 FILLER_12_943 ();
 sg13g2_decap_8 FILLER_12_950 ();
 sg13g2_decap_8 FILLER_12_957 ();
 sg13g2_decap_8 FILLER_12_964 ();
 sg13g2_decap_8 FILLER_12_971 ();
 sg13g2_decap_8 FILLER_12_978 ();
 sg13g2_decap_8 FILLER_12_985 ();
 sg13g2_decap_8 FILLER_12_992 ();
 sg13g2_decap_8 FILLER_12_999 ();
 sg13g2_decap_8 FILLER_12_1006 ();
 sg13g2_decap_8 FILLER_12_1013 ();
 sg13g2_decap_8 FILLER_12_1020 ();
 sg13g2_fill_2 FILLER_12_1027 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_fill_2 FILLER_13_67 ();
 sg13g2_fill_2 FILLER_13_96 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_decap_4 FILLER_13_141 ();
 sg13g2_fill_1 FILLER_13_145 ();
 sg13g2_decap_4 FILLER_13_165 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_decap_4 FILLER_13_230 ();
 sg13g2_fill_2 FILLER_13_234 ();
 sg13g2_fill_2 FILLER_13_243 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_260 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_decap_4 FILLER_13_288 ();
 sg13g2_fill_2 FILLER_13_315 ();
 sg13g2_fill_1 FILLER_13_317 ();
 sg13g2_decap_4 FILLER_13_326 ();
 sg13g2_fill_1 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_4 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_decap_8 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_13_868 ();
 sg13g2_decap_8 FILLER_13_875 ();
 sg13g2_decap_8 FILLER_13_882 ();
 sg13g2_decap_8 FILLER_13_889 ();
 sg13g2_decap_8 FILLER_13_896 ();
 sg13g2_decap_8 FILLER_13_903 ();
 sg13g2_decap_8 FILLER_13_910 ();
 sg13g2_decap_8 FILLER_13_917 ();
 sg13g2_decap_8 FILLER_13_924 ();
 sg13g2_decap_8 FILLER_13_931 ();
 sg13g2_decap_8 FILLER_13_938 ();
 sg13g2_decap_8 FILLER_13_945 ();
 sg13g2_decap_8 FILLER_13_952 ();
 sg13g2_decap_8 FILLER_13_959 ();
 sg13g2_decap_8 FILLER_13_966 ();
 sg13g2_decap_8 FILLER_13_973 ();
 sg13g2_decap_8 FILLER_13_980 ();
 sg13g2_decap_8 FILLER_13_987 ();
 sg13g2_decap_8 FILLER_13_994 ();
 sg13g2_decap_8 FILLER_13_1001 ();
 sg13g2_decap_8 FILLER_13_1008 ();
 sg13g2_decap_8 FILLER_13_1015 ();
 sg13g2_decap_8 FILLER_13_1022 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_fill_2 FILLER_14_53 ();
 sg13g2_fill_1 FILLER_14_55 ();
 sg13g2_fill_1 FILLER_14_83 ();
 sg13g2_fill_1 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_125 ();
 sg13g2_fill_2 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_143 ();
 sg13g2_decap_8 FILLER_14_171 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_fill_1 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_218 ();
 sg13g2_decap_4 FILLER_14_256 ();
 sg13g2_fill_2 FILLER_14_260 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_fill_1 FILLER_14_294 ();
 sg13g2_decap_4 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_327 ();
 sg13g2_decap_4 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_decap_8 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_14_436 ();
 sg13g2_decap_8 FILLER_14_443 ();
 sg13g2_decap_8 FILLER_14_450 ();
 sg13g2_decap_8 FILLER_14_457 ();
 sg13g2_decap_8 FILLER_14_464 ();
 sg13g2_decap_8 FILLER_14_471 ();
 sg13g2_decap_8 FILLER_14_478 ();
 sg13g2_decap_8 FILLER_14_485 ();
 sg13g2_decap_8 FILLER_14_492 ();
 sg13g2_decap_8 FILLER_14_499 ();
 sg13g2_decap_8 FILLER_14_506 ();
 sg13g2_decap_8 FILLER_14_513 ();
 sg13g2_decap_8 FILLER_14_520 ();
 sg13g2_decap_8 FILLER_14_527 ();
 sg13g2_decap_8 FILLER_14_534 ();
 sg13g2_decap_8 FILLER_14_541 ();
 sg13g2_decap_8 FILLER_14_548 ();
 sg13g2_decap_8 FILLER_14_555 ();
 sg13g2_decap_8 FILLER_14_562 ();
 sg13g2_decap_8 FILLER_14_569 ();
 sg13g2_decap_8 FILLER_14_576 ();
 sg13g2_decap_8 FILLER_14_583 ();
 sg13g2_decap_8 FILLER_14_590 ();
 sg13g2_decap_8 FILLER_14_597 ();
 sg13g2_decap_8 FILLER_14_604 ();
 sg13g2_decap_8 FILLER_14_611 ();
 sg13g2_decap_8 FILLER_14_618 ();
 sg13g2_decap_8 FILLER_14_625 ();
 sg13g2_decap_8 FILLER_14_632 ();
 sg13g2_decap_8 FILLER_14_639 ();
 sg13g2_decap_8 FILLER_14_646 ();
 sg13g2_decap_8 FILLER_14_653 ();
 sg13g2_decap_8 FILLER_14_660 ();
 sg13g2_decap_8 FILLER_14_667 ();
 sg13g2_decap_8 FILLER_14_674 ();
 sg13g2_decap_8 FILLER_14_681 ();
 sg13g2_decap_8 FILLER_14_688 ();
 sg13g2_decap_8 FILLER_14_695 ();
 sg13g2_decap_8 FILLER_14_702 ();
 sg13g2_decap_8 FILLER_14_709 ();
 sg13g2_decap_8 FILLER_14_716 ();
 sg13g2_decap_8 FILLER_14_723 ();
 sg13g2_decap_8 FILLER_14_730 ();
 sg13g2_decap_8 FILLER_14_737 ();
 sg13g2_decap_8 FILLER_14_744 ();
 sg13g2_decap_8 FILLER_14_751 ();
 sg13g2_decap_8 FILLER_14_758 ();
 sg13g2_decap_8 FILLER_14_765 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_decap_8 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_14_835 ();
 sg13g2_decap_8 FILLER_14_842 ();
 sg13g2_decap_8 FILLER_14_849 ();
 sg13g2_decap_8 FILLER_14_856 ();
 sg13g2_decap_8 FILLER_14_863 ();
 sg13g2_decap_8 FILLER_14_870 ();
 sg13g2_decap_8 FILLER_14_877 ();
 sg13g2_decap_8 FILLER_14_884 ();
 sg13g2_decap_8 FILLER_14_891 ();
 sg13g2_decap_8 FILLER_14_898 ();
 sg13g2_decap_8 FILLER_14_905 ();
 sg13g2_decap_8 FILLER_14_912 ();
 sg13g2_decap_8 FILLER_14_919 ();
 sg13g2_decap_8 FILLER_14_926 ();
 sg13g2_decap_8 FILLER_14_933 ();
 sg13g2_decap_8 FILLER_14_940 ();
 sg13g2_decap_8 FILLER_14_947 ();
 sg13g2_decap_8 FILLER_14_954 ();
 sg13g2_decap_8 FILLER_14_961 ();
 sg13g2_decap_8 FILLER_14_968 ();
 sg13g2_decap_8 FILLER_14_975 ();
 sg13g2_decap_8 FILLER_14_982 ();
 sg13g2_decap_8 FILLER_14_989 ();
 sg13g2_decap_8 FILLER_14_996 ();
 sg13g2_decap_8 FILLER_14_1003 ();
 sg13g2_decap_8 FILLER_14_1010 ();
 sg13g2_decap_8 FILLER_14_1017 ();
 sg13g2_decap_4 FILLER_14_1024 ();
 sg13g2_fill_1 FILLER_14_1028 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_fill_1 FILLER_15_36 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_1 FILLER_15_52 ();
 sg13g2_fill_1 FILLER_15_82 ();
 sg13g2_decap_4 FILLER_15_110 ();
 sg13g2_decap_4 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_decap_8 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_183 ();
 sg13g2_fill_1 FILLER_15_207 ();
 sg13g2_decap_4 FILLER_15_227 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_236 ();
 sg13g2_decap_8 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_fill_1 FILLER_15_325 ();
 sg13g2_decap_4 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_fill_2 FILLER_15_387 ();
 sg13g2_fill_1 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_473 ();
 sg13g2_decap_8 FILLER_15_480 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_494 ();
 sg13g2_decap_8 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_508 ();
 sg13g2_decap_8 FILLER_15_515 ();
 sg13g2_decap_8 FILLER_15_522 ();
 sg13g2_decap_8 FILLER_15_529 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_decap_8 FILLER_15_564 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_decap_8 FILLER_15_585 ();
 sg13g2_decap_8 FILLER_15_592 ();
 sg13g2_decap_8 FILLER_15_599 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_decap_8 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_697 ();
 sg13g2_decap_8 FILLER_15_704 ();
 sg13g2_decap_8 FILLER_15_711 ();
 sg13g2_decap_8 FILLER_15_718 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_decap_8 FILLER_15_739 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_decap_8 FILLER_15_753 ();
 sg13g2_decap_8 FILLER_15_760 ();
 sg13g2_decap_8 FILLER_15_767 ();
 sg13g2_decap_8 FILLER_15_774 ();
 sg13g2_decap_8 FILLER_15_781 ();
 sg13g2_decap_8 FILLER_15_788 ();
 sg13g2_decap_8 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_decap_8 FILLER_15_809 ();
 sg13g2_decap_8 FILLER_15_816 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_decap_8 FILLER_15_830 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_decap_8 FILLER_15_858 ();
 sg13g2_decap_8 FILLER_15_865 ();
 sg13g2_decap_8 FILLER_15_872 ();
 sg13g2_decap_8 FILLER_15_879 ();
 sg13g2_decap_8 FILLER_15_886 ();
 sg13g2_decap_8 FILLER_15_893 ();
 sg13g2_decap_8 FILLER_15_900 ();
 sg13g2_decap_8 FILLER_15_907 ();
 sg13g2_decap_8 FILLER_15_914 ();
 sg13g2_decap_8 FILLER_15_921 ();
 sg13g2_decap_8 FILLER_15_928 ();
 sg13g2_decap_8 FILLER_15_935 ();
 sg13g2_decap_8 FILLER_15_942 ();
 sg13g2_decap_8 FILLER_15_949 ();
 sg13g2_decap_8 FILLER_15_956 ();
 sg13g2_decap_8 FILLER_15_963 ();
 sg13g2_decap_8 FILLER_15_970 ();
 sg13g2_decap_8 FILLER_15_977 ();
 sg13g2_decap_8 FILLER_15_984 ();
 sg13g2_decap_8 FILLER_15_991 ();
 sg13g2_decap_8 FILLER_15_998 ();
 sg13g2_decap_8 FILLER_15_1005 ();
 sg13g2_decap_8 FILLER_15_1012 ();
 sg13g2_decap_8 FILLER_15_1019 ();
 sg13g2_fill_2 FILLER_15_1026 ();
 sg13g2_fill_1 FILLER_15_1028 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_8 FILLER_16_18 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_fill_2 FILLER_16_96 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_decap_4 FILLER_16_165 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_185 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_decap_4 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_255 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_2 FILLER_16_267 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_decap_4 FILLER_16_316 ();
 sg13g2_decap_4 FILLER_16_325 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_decap_4 FILLER_16_373 ();
 sg13g2_fill_1 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_decap_8 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_decap_8 FILLER_16_875 ();
 sg13g2_decap_8 FILLER_16_882 ();
 sg13g2_decap_8 FILLER_16_889 ();
 sg13g2_decap_8 FILLER_16_896 ();
 sg13g2_decap_8 FILLER_16_903 ();
 sg13g2_decap_8 FILLER_16_910 ();
 sg13g2_decap_8 FILLER_16_917 ();
 sg13g2_decap_8 FILLER_16_924 ();
 sg13g2_decap_8 FILLER_16_931 ();
 sg13g2_decap_8 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_945 ();
 sg13g2_decap_8 FILLER_16_952 ();
 sg13g2_decap_8 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_966 ();
 sg13g2_decap_8 FILLER_16_973 ();
 sg13g2_decap_8 FILLER_16_980 ();
 sg13g2_decap_8 FILLER_16_987 ();
 sg13g2_decap_8 FILLER_16_994 ();
 sg13g2_decap_8 FILLER_16_1001 ();
 sg13g2_decap_8 FILLER_16_1008 ();
 sg13g2_decap_8 FILLER_16_1015 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_32 ();
 sg13g2_fill_1 FILLER_17_83 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_236 ();
 sg13g2_decap_8 FILLER_17_243 ();
 sg13g2_decap_8 FILLER_17_250 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_decap_4 FILLER_17_268 ();
 sg13g2_fill_1 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_4 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_8 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_17_431 ();
 sg13g2_decap_8 FILLER_17_438 ();
 sg13g2_decap_8 FILLER_17_445 ();
 sg13g2_decap_8 FILLER_17_452 ();
 sg13g2_decap_8 FILLER_17_459 ();
 sg13g2_decap_8 FILLER_17_466 ();
 sg13g2_decap_8 FILLER_17_473 ();
 sg13g2_decap_8 FILLER_17_480 ();
 sg13g2_decap_8 FILLER_17_487 ();
 sg13g2_decap_8 FILLER_17_494 ();
 sg13g2_decap_8 FILLER_17_501 ();
 sg13g2_decap_8 FILLER_17_508 ();
 sg13g2_decap_8 FILLER_17_515 ();
 sg13g2_decap_8 FILLER_17_522 ();
 sg13g2_decap_8 FILLER_17_529 ();
 sg13g2_decap_8 FILLER_17_536 ();
 sg13g2_decap_8 FILLER_17_543 ();
 sg13g2_decap_8 FILLER_17_550 ();
 sg13g2_decap_8 FILLER_17_557 ();
 sg13g2_decap_8 FILLER_17_564 ();
 sg13g2_decap_8 FILLER_17_571 ();
 sg13g2_decap_8 FILLER_17_578 ();
 sg13g2_decap_8 FILLER_17_585 ();
 sg13g2_decap_8 FILLER_17_592 ();
 sg13g2_decap_8 FILLER_17_599 ();
 sg13g2_decap_8 FILLER_17_606 ();
 sg13g2_decap_8 FILLER_17_613 ();
 sg13g2_decap_8 FILLER_17_620 ();
 sg13g2_decap_8 FILLER_17_627 ();
 sg13g2_decap_8 FILLER_17_634 ();
 sg13g2_decap_8 FILLER_17_641 ();
 sg13g2_decap_8 FILLER_17_648 ();
 sg13g2_decap_8 FILLER_17_655 ();
 sg13g2_decap_8 FILLER_17_662 ();
 sg13g2_decap_8 FILLER_17_669 ();
 sg13g2_decap_8 FILLER_17_676 ();
 sg13g2_decap_8 FILLER_17_683 ();
 sg13g2_decap_8 FILLER_17_690 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_decap_8 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_711 ();
 sg13g2_decap_8 FILLER_17_718 ();
 sg13g2_decap_8 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_732 ();
 sg13g2_decap_8 FILLER_17_739 ();
 sg13g2_decap_8 FILLER_17_746 ();
 sg13g2_decap_8 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_decap_8 FILLER_17_774 ();
 sg13g2_decap_8 FILLER_17_781 ();
 sg13g2_decap_8 FILLER_17_788 ();
 sg13g2_decap_8 FILLER_17_795 ();
 sg13g2_decap_8 FILLER_17_802 ();
 sg13g2_decap_8 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_decap_8 FILLER_17_830 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_decap_8 FILLER_17_844 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_decap_8 FILLER_17_858 ();
 sg13g2_decap_8 FILLER_17_865 ();
 sg13g2_decap_8 FILLER_17_872 ();
 sg13g2_decap_8 FILLER_17_879 ();
 sg13g2_decap_8 FILLER_17_886 ();
 sg13g2_decap_8 FILLER_17_893 ();
 sg13g2_decap_8 FILLER_17_900 ();
 sg13g2_decap_8 FILLER_17_907 ();
 sg13g2_decap_8 FILLER_17_914 ();
 sg13g2_decap_8 FILLER_17_921 ();
 sg13g2_decap_8 FILLER_17_928 ();
 sg13g2_decap_8 FILLER_17_935 ();
 sg13g2_decap_8 FILLER_17_942 ();
 sg13g2_decap_8 FILLER_17_949 ();
 sg13g2_decap_8 FILLER_17_956 ();
 sg13g2_decap_8 FILLER_17_963 ();
 sg13g2_decap_8 FILLER_17_970 ();
 sg13g2_decap_8 FILLER_17_977 ();
 sg13g2_decap_8 FILLER_17_984 ();
 sg13g2_decap_8 FILLER_17_991 ();
 sg13g2_decap_8 FILLER_17_998 ();
 sg13g2_decap_8 FILLER_17_1005 ();
 sg13g2_decap_8 FILLER_17_1012 ();
 sg13g2_decap_8 FILLER_17_1019 ();
 sg13g2_fill_2 FILLER_17_1026 ();
 sg13g2_fill_1 FILLER_17_1028 ();
 sg13g2_fill_1 FILLER_18_8 ();
 sg13g2_decap_8 FILLER_18_13 ();
 sg13g2_decap_4 FILLER_18_20 ();
 sg13g2_decap_4 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_103 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_4 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_134 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_decap_4 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_4 FILLER_18_361 ();
 sg13g2_decap_4 FILLER_18_376 ();
 sg13g2_fill_2 FILLER_18_393 ();
 sg13g2_fill_1 FILLER_18_395 ();
 sg13g2_fill_1 FILLER_18_400 ();
 sg13g2_decap_8 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_18_436 ();
 sg13g2_decap_8 FILLER_18_443 ();
 sg13g2_decap_8 FILLER_18_450 ();
 sg13g2_decap_8 FILLER_18_457 ();
 sg13g2_decap_8 FILLER_18_464 ();
 sg13g2_decap_8 FILLER_18_471 ();
 sg13g2_decap_8 FILLER_18_478 ();
 sg13g2_decap_8 FILLER_18_485 ();
 sg13g2_decap_8 FILLER_18_492 ();
 sg13g2_decap_8 FILLER_18_499 ();
 sg13g2_decap_8 FILLER_18_506 ();
 sg13g2_decap_8 FILLER_18_513 ();
 sg13g2_decap_8 FILLER_18_520 ();
 sg13g2_decap_8 FILLER_18_527 ();
 sg13g2_decap_8 FILLER_18_534 ();
 sg13g2_decap_8 FILLER_18_541 ();
 sg13g2_decap_8 FILLER_18_548 ();
 sg13g2_decap_8 FILLER_18_555 ();
 sg13g2_decap_8 FILLER_18_562 ();
 sg13g2_decap_8 FILLER_18_569 ();
 sg13g2_decap_8 FILLER_18_576 ();
 sg13g2_decap_8 FILLER_18_583 ();
 sg13g2_decap_8 FILLER_18_590 ();
 sg13g2_decap_8 FILLER_18_597 ();
 sg13g2_decap_8 FILLER_18_604 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_decap_8 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_625 ();
 sg13g2_decap_8 FILLER_18_632 ();
 sg13g2_decap_8 FILLER_18_639 ();
 sg13g2_decap_8 FILLER_18_646 ();
 sg13g2_decap_8 FILLER_18_653 ();
 sg13g2_decap_8 FILLER_18_660 ();
 sg13g2_decap_8 FILLER_18_667 ();
 sg13g2_decap_8 FILLER_18_674 ();
 sg13g2_decap_8 FILLER_18_681 ();
 sg13g2_decap_8 FILLER_18_688 ();
 sg13g2_decap_8 FILLER_18_695 ();
 sg13g2_decap_8 FILLER_18_702 ();
 sg13g2_decap_8 FILLER_18_709 ();
 sg13g2_decap_8 FILLER_18_716 ();
 sg13g2_decap_8 FILLER_18_723 ();
 sg13g2_decap_8 FILLER_18_730 ();
 sg13g2_decap_8 FILLER_18_737 ();
 sg13g2_decap_8 FILLER_18_744 ();
 sg13g2_decap_8 FILLER_18_751 ();
 sg13g2_decap_8 FILLER_18_758 ();
 sg13g2_decap_8 FILLER_18_765 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_8 FILLER_18_779 ();
 sg13g2_decap_8 FILLER_18_786 ();
 sg13g2_decap_8 FILLER_18_793 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_decap_8 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_842 ();
 sg13g2_decap_8 FILLER_18_849 ();
 sg13g2_decap_8 FILLER_18_856 ();
 sg13g2_decap_8 FILLER_18_863 ();
 sg13g2_decap_8 FILLER_18_870 ();
 sg13g2_decap_8 FILLER_18_877 ();
 sg13g2_decap_8 FILLER_18_884 ();
 sg13g2_decap_8 FILLER_18_891 ();
 sg13g2_decap_8 FILLER_18_898 ();
 sg13g2_decap_8 FILLER_18_905 ();
 sg13g2_decap_8 FILLER_18_912 ();
 sg13g2_decap_8 FILLER_18_919 ();
 sg13g2_decap_8 FILLER_18_926 ();
 sg13g2_decap_8 FILLER_18_933 ();
 sg13g2_decap_8 FILLER_18_940 ();
 sg13g2_decap_8 FILLER_18_947 ();
 sg13g2_decap_8 FILLER_18_954 ();
 sg13g2_decap_8 FILLER_18_961 ();
 sg13g2_decap_8 FILLER_18_968 ();
 sg13g2_decap_8 FILLER_18_975 ();
 sg13g2_decap_8 FILLER_18_982 ();
 sg13g2_decap_8 FILLER_18_989 ();
 sg13g2_decap_8 FILLER_18_996 ();
 sg13g2_decap_8 FILLER_18_1003 ();
 sg13g2_decap_8 FILLER_18_1010 ();
 sg13g2_decap_8 FILLER_18_1017 ();
 sg13g2_decap_4 FILLER_18_1024 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_31 ();
 sg13g2_fill_1 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_117 ();
 sg13g2_decap_4 FILLER_19_124 ();
 sg13g2_decap_8 FILLER_19_173 ();
 sg13g2_decap_8 FILLER_19_180 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_236 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_fill_2 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_250 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_4 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_308 ();
 sg13g2_fill_1 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_fill_2 FILLER_19_338 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_360 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_418 ();
 sg13g2_decap_8 FILLER_19_425 ();
 sg13g2_decap_8 FILLER_19_432 ();
 sg13g2_decap_8 FILLER_19_439 ();
 sg13g2_decap_8 FILLER_19_446 ();
 sg13g2_decap_8 FILLER_19_453 ();
 sg13g2_decap_8 FILLER_19_460 ();
 sg13g2_decap_8 FILLER_19_467 ();
 sg13g2_decap_8 FILLER_19_474 ();
 sg13g2_decap_8 FILLER_19_481 ();
 sg13g2_decap_8 FILLER_19_488 ();
 sg13g2_decap_8 FILLER_19_495 ();
 sg13g2_decap_8 FILLER_19_502 ();
 sg13g2_decap_8 FILLER_19_509 ();
 sg13g2_decap_8 FILLER_19_516 ();
 sg13g2_decap_8 FILLER_19_523 ();
 sg13g2_decap_8 FILLER_19_530 ();
 sg13g2_decap_8 FILLER_19_537 ();
 sg13g2_decap_8 FILLER_19_544 ();
 sg13g2_decap_8 FILLER_19_551 ();
 sg13g2_decap_8 FILLER_19_558 ();
 sg13g2_decap_8 FILLER_19_565 ();
 sg13g2_decap_8 FILLER_19_572 ();
 sg13g2_decap_8 FILLER_19_579 ();
 sg13g2_decap_8 FILLER_19_586 ();
 sg13g2_decap_8 FILLER_19_593 ();
 sg13g2_decap_8 FILLER_19_600 ();
 sg13g2_decap_8 FILLER_19_607 ();
 sg13g2_decap_8 FILLER_19_614 ();
 sg13g2_decap_8 FILLER_19_621 ();
 sg13g2_decap_8 FILLER_19_628 ();
 sg13g2_decap_8 FILLER_19_635 ();
 sg13g2_decap_8 FILLER_19_642 ();
 sg13g2_decap_8 FILLER_19_649 ();
 sg13g2_decap_8 FILLER_19_656 ();
 sg13g2_decap_8 FILLER_19_663 ();
 sg13g2_decap_8 FILLER_19_670 ();
 sg13g2_decap_8 FILLER_19_677 ();
 sg13g2_decap_8 FILLER_19_684 ();
 sg13g2_decap_8 FILLER_19_691 ();
 sg13g2_decap_8 FILLER_19_698 ();
 sg13g2_decap_8 FILLER_19_705 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_719 ();
 sg13g2_decap_8 FILLER_19_726 ();
 sg13g2_decap_8 FILLER_19_733 ();
 sg13g2_decap_8 FILLER_19_740 ();
 sg13g2_decap_8 FILLER_19_747 ();
 sg13g2_decap_8 FILLER_19_754 ();
 sg13g2_decap_8 FILLER_19_761 ();
 sg13g2_decap_8 FILLER_19_768 ();
 sg13g2_decap_8 FILLER_19_775 ();
 sg13g2_decap_8 FILLER_19_782 ();
 sg13g2_decap_8 FILLER_19_789 ();
 sg13g2_decap_8 FILLER_19_796 ();
 sg13g2_decap_8 FILLER_19_803 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_decap_8 FILLER_19_824 ();
 sg13g2_decap_8 FILLER_19_831 ();
 sg13g2_decap_8 FILLER_19_838 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_decap_8 FILLER_19_859 ();
 sg13g2_decap_8 FILLER_19_866 ();
 sg13g2_decap_8 FILLER_19_873 ();
 sg13g2_decap_8 FILLER_19_880 ();
 sg13g2_decap_8 FILLER_19_887 ();
 sg13g2_decap_8 FILLER_19_894 ();
 sg13g2_decap_8 FILLER_19_901 ();
 sg13g2_decap_8 FILLER_19_908 ();
 sg13g2_decap_8 FILLER_19_915 ();
 sg13g2_decap_8 FILLER_19_922 ();
 sg13g2_decap_8 FILLER_19_929 ();
 sg13g2_decap_8 FILLER_19_936 ();
 sg13g2_decap_8 FILLER_19_943 ();
 sg13g2_decap_8 FILLER_19_950 ();
 sg13g2_decap_8 FILLER_19_957 ();
 sg13g2_decap_8 FILLER_19_964 ();
 sg13g2_decap_8 FILLER_19_971 ();
 sg13g2_decap_8 FILLER_19_978 ();
 sg13g2_decap_8 FILLER_19_985 ();
 sg13g2_decap_8 FILLER_19_992 ();
 sg13g2_decap_8 FILLER_19_999 ();
 sg13g2_decap_8 FILLER_19_1006 ();
 sg13g2_decap_8 FILLER_19_1013 ();
 sg13g2_decap_8 FILLER_19_1020 ();
 sg13g2_fill_2 FILLER_19_1027 ();
 sg13g2_decap_4 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_12 ();
 sg13g2_decap_4 FILLER_20_19 ();
 sg13g2_fill_2 FILLER_20_23 ();
 sg13g2_fill_1 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_65 ();
 sg13g2_fill_1 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_118 ();
 sg13g2_fill_2 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_176 ();
 sg13g2_decap_4 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_220 ();
 sg13g2_decap_8 FILLER_20_254 ();
 sg13g2_decap_4 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_294 ();
 sg13g2_decap_4 FILLER_20_300 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_352 ();
 sg13g2_fill_2 FILLER_20_376 ();
 sg13g2_fill_2 FILLER_20_387 ();
 sg13g2_fill_2 FILLER_20_396 ();
 sg13g2_fill_1 FILLER_20_398 ();
 sg13g2_decap_8 FILLER_20_426 ();
 sg13g2_decap_8 FILLER_20_433 ();
 sg13g2_decap_8 FILLER_20_440 ();
 sg13g2_decap_8 FILLER_20_447 ();
 sg13g2_decap_8 FILLER_20_454 ();
 sg13g2_decap_8 FILLER_20_461 ();
 sg13g2_decap_8 FILLER_20_468 ();
 sg13g2_decap_8 FILLER_20_475 ();
 sg13g2_decap_8 FILLER_20_482 ();
 sg13g2_decap_8 FILLER_20_489 ();
 sg13g2_decap_8 FILLER_20_496 ();
 sg13g2_decap_8 FILLER_20_503 ();
 sg13g2_decap_8 FILLER_20_510 ();
 sg13g2_decap_8 FILLER_20_517 ();
 sg13g2_decap_8 FILLER_20_524 ();
 sg13g2_decap_8 FILLER_20_531 ();
 sg13g2_decap_8 FILLER_20_538 ();
 sg13g2_decap_8 FILLER_20_545 ();
 sg13g2_decap_8 FILLER_20_552 ();
 sg13g2_decap_8 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_566 ();
 sg13g2_decap_8 FILLER_20_573 ();
 sg13g2_decap_8 FILLER_20_580 ();
 sg13g2_decap_8 FILLER_20_587 ();
 sg13g2_decap_8 FILLER_20_594 ();
 sg13g2_decap_8 FILLER_20_601 ();
 sg13g2_decap_8 FILLER_20_608 ();
 sg13g2_decap_8 FILLER_20_615 ();
 sg13g2_decap_8 FILLER_20_622 ();
 sg13g2_decap_8 FILLER_20_629 ();
 sg13g2_decap_8 FILLER_20_636 ();
 sg13g2_decap_8 FILLER_20_643 ();
 sg13g2_decap_8 FILLER_20_650 ();
 sg13g2_decap_8 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_664 ();
 sg13g2_decap_8 FILLER_20_671 ();
 sg13g2_decap_8 FILLER_20_678 ();
 sg13g2_decap_8 FILLER_20_685 ();
 sg13g2_decap_8 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_699 ();
 sg13g2_decap_8 FILLER_20_706 ();
 sg13g2_decap_8 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_720 ();
 sg13g2_decap_8 FILLER_20_727 ();
 sg13g2_decap_8 FILLER_20_734 ();
 sg13g2_decap_8 FILLER_20_741 ();
 sg13g2_decap_8 FILLER_20_748 ();
 sg13g2_decap_8 FILLER_20_755 ();
 sg13g2_decap_8 FILLER_20_762 ();
 sg13g2_decap_8 FILLER_20_769 ();
 sg13g2_decap_8 FILLER_20_776 ();
 sg13g2_decap_8 FILLER_20_783 ();
 sg13g2_decap_8 FILLER_20_790 ();
 sg13g2_decap_8 FILLER_20_797 ();
 sg13g2_decap_8 FILLER_20_804 ();
 sg13g2_decap_8 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_818 ();
 sg13g2_decap_8 FILLER_20_825 ();
 sg13g2_decap_8 FILLER_20_832 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_decap_8 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_20_867 ();
 sg13g2_decap_8 FILLER_20_874 ();
 sg13g2_decap_8 FILLER_20_881 ();
 sg13g2_decap_8 FILLER_20_888 ();
 sg13g2_decap_8 FILLER_20_895 ();
 sg13g2_decap_8 FILLER_20_902 ();
 sg13g2_decap_8 FILLER_20_909 ();
 sg13g2_decap_8 FILLER_20_916 ();
 sg13g2_decap_8 FILLER_20_923 ();
 sg13g2_decap_8 FILLER_20_930 ();
 sg13g2_decap_8 FILLER_20_937 ();
 sg13g2_decap_8 FILLER_20_944 ();
 sg13g2_decap_8 FILLER_20_951 ();
 sg13g2_decap_8 FILLER_20_958 ();
 sg13g2_decap_8 FILLER_20_965 ();
 sg13g2_decap_8 FILLER_20_972 ();
 sg13g2_decap_8 FILLER_20_979 ();
 sg13g2_decap_8 FILLER_20_986 ();
 sg13g2_decap_8 FILLER_20_993 ();
 sg13g2_decap_8 FILLER_20_1000 ();
 sg13g2_decap_8 FILLER_20_1007 ();
 sg13g2_decap_8 FILLER_20_1014 ();
 sg13g2_decap_8 FILLER_20_1021 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_fill_2 FILLER_21_25 ();
 sg13g2_fill_2 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_4 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_2 FILLER_21_100 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_2 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_193 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_4 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_261 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_291 ();
 sg13g2_decap_4 FILLER_21_313 ();
 sg13g2_decap_4 FILLER_21_361 ();
 sg13g2_fill_2 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_437 ();
 sg13g2_decap_8 FILLER_21_444 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_decap_8 FILLER_21_458 ();
 sg13g2_decap_8 FILLER_21_465 ();
 sg13g2_decap_8 FILLER_21_472 ();
 sg13g2_decap_8 FILLER_21_479 ();
 sg13g2_decap_8 FILLER_21_486 ();
 sg13g2_decap_8 FILLER_21_493 ();
 sg13g2_decap_8 FILLER_21_500 ();
 sg13g2_decap_8 FILLER_21_507 ();
 sg13g2_decap_8 FILLER_21_514 ();
 sg13g2_decap_8 FILLER_21_521 ();
 sg13g2_decap_8 FILLER_21_528 ();
 sg13g2_decap_8 FILLER_21_535 ();
 sg13g2_decap_8 FILLER_21_542 ();
 sg13g2_decap_8 FILLER_21_549 ();
 sg13g2_decap_8 FILLER_21_556 ();
 sg13g2_decap_8 FILLER_21_563 ();
 sg13g2_decap_8 FILLER_21_570 ();
 sg13g2_decap_8 FILLER_21_577 ();
 sg13g2_decap_8 FILLER_21_584 ();
 sg13g2_decap_8 FILLER_21_591 ();
 sg13g2_decap_8 FILLER_21_598 ();
 sg13g2_decap_8 FILLER_21_605 ();
 sg13g2_decap_8 FILLER_21_612 ();
 sg13g2_decap_8 FILLER_21_619 ();
 sg13g2_decap_8 FILLER_21_626 ();
 sg13g2_decap_8 FILLER_21_633 ();
 sg13g2_decap_8 FILLER_21_640 ();
 sg13g2_decap_8 FILLER_21_647 ();
 sg13g2_decap_8 FILLER_21_654 ();
 sg13g2_decap_8 FILLER_21_661 ();
 sg13g2_decap_8 FILLER_21_668 ();
 sg13g2_decap_8 FILLER_21_675 ();
 sg13g2_decap_8 FILLER_21_682 ();
 sg13g2_decap_8 FILLER_21_689 ();
 sg13g2_decap_8 FILLER_21_696 ();
 sg13g2_decap_8 FILLER_21_703 ();
 sg13g2_decap_8 FILLER_21_710 ();
 sg13g2_decap_8 FILLER_21_717 ();
 sg13g2_decap_8 FILLER_21_724 ();
 sg13g2_decap_8 FILLER_21_731 ();
 sg13g2_decap_8 FILLER_21_738 ();
 sg13g2_decap_8 FILLER_21_745 ();
 sg13g2_decap_8 FILLER_21_752 ();
 sg13g2_decap_8 FILLER_21_759 ();
 sg13g2_decap_8 FILLER_21_766 ();
 sg13g2_decap_8 FILLER_21_773 ();
 sg13g2_decap_8 FILLER_21_780 ();
 sg13g2_decap_8 FILLER_21_787 ();
 sg13g2_decap_8 FILLER_21_794 ();
 sg13g2_decap_8 FILLER_21_801 ();
 sg13g2_decap_8 FILLER_21_808 ();
 sg13g2_decap_8 FILLER_21_815 ();
 sg13g2_decap_8 FILLER_21_822 ();
 sg13g2_decap_8 FILLER_21_829 ();
 sg13g2_decap_8 FILLER_21_836 ();
 sg13g2_decap_8 FILLER_21_843 ();
 sg13g2_decap_8 FILLER_21_850 ();
 sg13g2_decap_8 FILLER_21_857 ();
 sg13g2_decap_8 FILLER_21_864 ();
 sg13g2_decap_8 FILLER_21_871 ();
 sg13g2_decap_8 FILLER_21_878 ();
 sg13g2_decap_8 FILLER_21_885 ();
 sg13g2_decap_8 FILLER_21_892 ();
 sg13g2_decap_8 FILLER_21_899 ();
 sg13g2_decap_8 FILLER_21_906 ();
 sg13g2_decap_8 FILLER_21_913 ();
 sg13g2_decap_8 FILLER_21_920 ();
 sg13g2_decap_8 FILLER_21_927 ();
 sg13g2_decap_8 FILLER_21_934 ();
 sg13g2_decap_8 FILLER_21_941 ();
 sg13g2_decap_8 FILLER_21_948 ();
 sg13g2_decap_8 FILLER_21_955 ();
 sg13g2_decap_8 FILLER_21_962 ();
 sg13g2_decap_8 FILLER_21_969 ();
 sg13g2_decap_8 FILLER_21_976 ();
 sg13g2_decap_8 FILLER_21_983 ();
 sg13g2_decap_8 FILLER_21_990 ();
 sg13g2_decap_8 FILLER_21_997 ();
 sg13g2_decap_8 FILLER_21_1004 ();
 sg13g2_decap_8 FILLER_21_1011 ();
 sg13g2_decap_8 FILLER_21_1018 ();
 sg13g2_decap_4 FILLER_21_1025 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_1 FILLER_22_38 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_fill_2 FILLER_22_113 ();
 sg13g2_decap_4 FILLER_22_152 ();
 sg13g2_fill_2 FILLER_22_156 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_decap_4 FILLER_22_343 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_425 ();
 sg13g2_decap_8 FILLER_22_432 ();
 sg13g2_decap_8 FILLER_22_439 ();
 sg13g2_decap_8 FILLER_22_446 ();
 sg13g2_decap_8 FILLER_22_453 ();
 sg13g2_decap_8 FILLER_22_460 ();
 sg13g2_decap_8 FILLER_22_467 ();
 sg13g2_decap_8 FILLER_22_474 ();
 sg13g2_decap_8 FILLER_22_481 ();
 sg13g2_decap_8 FILLER_22_488 ();
 sg13g2_decap_8 FILLER_22_495 ();
 sg13g2_decap_8 FILLER_22_502 ();
 sg13g2_decap_8 FILLER_22_509 ();
 sg13g2_decap_8 FILLER_22_516 ();
 sg13g2_decap_8 FILLER_22_523 ();
 sg13g2_decap_8 FILLER_22_530 ();
 sg13g2_decap_8 FILLER_22_537 ();
 sg13g2_decap_8 FILLER_22_544 ();
 sg13g2_decap_8 FILLER_22_551 ();
 sg13g2_decap_8 FILLER_22_558 ();
 sg13g2_decap_8 FILLER_22_565 ();
 sg13g2_decap_8 FILLER_22_572 ();
 sg13g2_decap_8 FILLER_22_579 ();
 sg13g2_decap_8 FILLER_22_586 ();
 sg13g2_decap_8 FILLER_22_593 ();
 sg13g2_decap_8 FILLER_22_600 ();
 sg13g2_decap_8 FILLER_22_607 ();
 sg13g2_decap_8 FILLER_22_614 ();
 sg13g2_decap_8 FILLER_22_621 ();
 sg13g2_decap_8 FILLER_22_628 ();
 sg13g2_decap_8 FILLER_22_635 ();
 sg13g2_decap_8 FILLER_22_642 ();
 sg13g2_decap_8 FILLER_22_649 ();
 sg13g2_decap_8 FILLER_22_656 ();
 sg13g2_decap_8 FILLER_22_663 ();
 sg13g2_decap_8 FILLER_22_670 ();
 sg13g2_decap_8 FILLER_22_677 ();
 sg13g2_decap_8 FILLER_22_684 ();
 sg13g2_decap_8 FILLER_22_691 ();
 sg13g2_decap_8 FILLER_22_698 ();
 sg13g2_decap_8 FILLER_22_705 ();
 sg13g2_decap_8 FILLER_22_712 ();
 sg13g2_decap_8 FILLER_22_719 ();
 sg13g2_decap_8 FILLER_22_726 ();
 sg13g2_decap_8 FILLER_22_733 ();
 sg13g2_decap_8 FILLER_22_740 ();
 sg13g2_decap_8 FILLER_22_747 ();
 sg13g2_decap_8 FILLER_22_754 ();
 sg13g2_decap_8 FILLER_22_761 ();
 sg13g2_decap_8 FILLER_22_768 ();
 sg13g2_decap_8 FILLER_22_775 ();
 sg13g2_decap_8 FILLER_22_782 ();
 sg13g2_decap_8 FILLER_22_789 ();
 sg13g2_decap_8 FILLER_22_796 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_decap_8 FILLER_22_810 ();
 sg13g2_decap_8 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_decap_8 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_838 ();
 sg13g2_decap_8 FILLER_22_845 ();
 sg13g2_decap_8 FILLER_22_852 ();
 sg13g2_decap_8 FILLER_22_859 ();
 sg13g2_decap_8 FILLER_22_866 ();
 sg13g2_decap_8 FILLER_22_873 ();
 sg13g2_decap_8 FILLER_22_880 ();
 sg13g2_decap_8 FILLER_22_887 ();
 sg13g2_decap_8 FILLER_22_894 ();
 sg13g2_decap_8 FILLER_22_901 ();
 sg13g2_decap_8 FILLER_22_908 ();
 sg13g2_decap_8 FILLER_22_915 ();
 sg13g2_decap_8 FILLER_22_922 ();
 sg13g2_decap_8 FILLER_22_929 ();
 sg13g2_decap_8 FILLER_22_936 ();
 sg13g2_decap_8 FILLER_22_943 ();
 sg13g2_decap_8 FILLER_22_950 ();
 sg13g2_decap_8 FILLER_22_957 ();
 sg13g2_decap_8 FILLER_22_964 ();
 sg13g2_decap_8 FILLER_22_971 ();
 sg13g2_decap_8 FILLER_22_978 ();
 sg13g2_decap_8 FILLER_22_985 ();
 sg13g2_decap_8 FILLER_22_992 ();
 sg13g2_decap_8 FILLER_22_999 ();
 sg13g2_decap_8 FILLER_22_1006 ();
 sg13g2_decap_8 FILLER_22_1013 ();
 sg13g2_decap_8 FILLER_22_1020 ();
 sg13g2_fill_2 FILLER_22_1027 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_6 ();
 sg13g2_fill_2 FILLER_23_48 ();
 sg13g2_fill_1 FILLER_23_50 ();
 sg13g2_decap_8 FILLER_23_78 ();
 sg13g2_decap_4 FILLER_23_85 ();
 sg13g2_fill_2 FILLER_23_89 ();
 sg13g2_decap_4 FILLER_23_95 ();
 sg13g2_fill_1 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_105 ();
 sg13g2_decap_4 FILLER_23_145 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_180 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_231 ();
 sg13g2_fill_1 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_342 ();
 sg13g2_fill_2 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_decap_8 FILLER_23_875 ();
 sg13g2_decap_8 FILLER_23_882 ();
 sg13g2_decap_8 FILLER_23_889 ();
 sg13g2_decap_8 FILLER_23_896 ();
 sg13g2_decap_8 FILLER_23_903 ();
 sg13g2_decap_8 FILLER_23_910 ();
 sg13g2_decap_8 FILLER_23_917 ();
 sg13g2_decap_8 FILLER_23_924 ();
 sg13g2_decap_8 FILLER_23_931 ();
 sg13g2_decap_8 FILLER_23_938 ();
 sg13g2_decap_8 FILLER_23_945 ();
 sg13g2_decap_8 FILLER_23_952 ();
 sg13g2_decap_8 FILLER_23_959 ();
 sg13g2_decap_8 FILLER_23_966 ();
 sg13g2_decap_8 FILLER_23_973 ();
 sg13g2_decap_8 FILLER_23_980 ();
 sg13g2_decap_8 FILLER_23_987 ();
 sg13g2_decap_8 FILLER_23_994 ();
 sg13g2_decap_8 FILLER_23_1001 ();
 sg13g2_decap_8 FILLER_23_1008 ();
 sg13g2_decap_8 FILLER_23_1015 ();
 sg13g2_decap_8 FILLER_23_1022 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_11 ();
 sg13g2_fill_1 FILLER_24_13 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_4 FILLER_24_25 ();
 sg13g2_fill_1 FILLER_24_29 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_4 FILLER_24_95 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_113 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_fill_2 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_2 FILLER_24_343 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_419 ();
 sg13g2_decap_8 FILLER_24_426 ();
 sg13g2_decap_8 FILLER_24_433 ();
 sg13g2_decap_8 FILLER_24_440 ();
 sg13g2_decap_8 FILLER_24_447 ();
 sg13g2_decap_8 FILLER_24_454 ();
 sg13g2_decap_8 FILLER_24_461 ();
 sg13g2_decap_8 FILLER_24_468 ();
 sg13g2_decap_8 FILLER_24_475 ();
 sg13g2_decap_8 FILLER_24_482 ();
 sg13g2_decap_8 FILLER_24_489 ();
 sg13g2_decap_8 FILLER_24_496 ();
 sg13g2_decap_8 FILLER_24_503 ();
 sg13g2_decap_8 FILLER_24_510 ();
 sg13g2_decap_8 FILLER_24_517 ();
 sg13g2_decap_8 FILLER_24_524 ();
 sg13g2_decap_8 FILLER_24_531 ();
 sg13g2_decap_8 FILLER_24_538 ();
 sg13g2_decap_8 FILLER_24_545 ();
 sg13g2_decap_8 FILLER_24_552 ();
 sg13g2_decap_8 FILLER_24_559 ();
 sg13g2_decap_8 FILLER_24_566 ();
 sg13g2_decap_8 FILLER_24_573 ();
 sg13g2_decap_8 FILLER_24_580 ();
 sg13g2_decap_8 FILLER_24_587 ();
 sg13g2_decap_8 FILLER_24_594 ();
 sg13g2_decap_8 FILLER_24_601 ();
 sg13g2_decap_8 FILLER_24_608 ();
 sg13g2_decap_8 FILLER_24_615 ();
 sg13g2_decap_8 FILLER_24_622 ();
 sg13g2_decap_8 FILLER_24_629 ();
 sg13g2_decap_8 FILLER_24_636 ();
 sg13g2_decap_8 FILLER_24_643 ();
 sg13g2_decap_8 FILLER_24_650 ();
 sg13g2_decap_8 FILLER_24_657 ();
 sg13g2_decap_8 FILLER_24_664 ();
 sg13g2_decap_8 FILLER_24_671 ();
 sg13g2_decap_8 FILLER_24_678 ();
 sg13g2_decap_8 FILLER_24_685 ();
 sg13g2_decap_8 FILLER_24_692 ();
 sg13g2_decap_8 FILLER_24_699 ();
 sg13g2_decap_8 FILLER_24_706 ();
 sg13g2_decap_8 FILLER_24_713 ();
 sg13g2_decap_8 FILLER_24_720 ();
 sg13g2_decap_8 FILLER_24_727 ();
 sg13g2_decap_8 FILLER_24_734 ();
 sg13g2_decap_8 FILLER_24_741 ();
 sg13g2_decap_8 FILLER_24_748 ();
 sg13g2_decap_8 FILLER_24_755 ();
 sg13g2_decap_8 FILLER_24_762 ();
 sg13g2_decap_8 FILLER_24_769 ();
 sg13g2_decap_8 FILLER_24_776 ();
 sg13g2_decap_8 FILLER_24_783 ();
 sg13g2_decap_8 FILLER_24_790 ();
 sg13g2_decap_8 FILLER_24_797 ();
 sg13g2_decap_8 FILLER_24_804 ();
 sg13g2_decap_8 FILLER_24_811 ();
 sg13g2_decap_8 FILLER_24_818 ();
 sg13g2_decap_8 FILLER_24_825 ();
 sg13g2_decap_8 FILLER_24_832 ();
 sg13g2_decap_8 FILLER_24_839 ();
 sg13g2_decap_8 FILLER_24_846 ();
 sg13g2_decap_8 FILLER_24_853 ();
 sg13g2_decap_8 FILLER_24_860 ();
 sg13g2_decap_8 FILLER_24_867 ();
 sg13g2_decap_8 FILLER_24_874 ();
 sg13g2_decap_8 FILLER_24_881 ();
 sg13g2_decap_8 FILLER_24_888 ();
 sg13g2_decap_8 FILLER_24_895 ();
 sg13g2_decap_8 FILLER_24_902 ();
 sg13g2_decap_8 FILLER_24_909 ();
 sg13g2_decap_8 FILLER_24_916 ();
 sg13g2_decap_8 FILLER_24_923 ();
 sg13g2_decap_8 FILLER_24_930 ();
 sg13g2_decap_8 FILLER_24_937 ();
 sg13g2_decap_8 FILLER_24_944 ();
 sg13g2_decap_8 FILLER_24_951 ();
 sg13g2_decap_8 FILLER_24_958 ();
 sg13g2_decap_8 FILLER_24_965 ();
 sg13g2_decap_8 FILLER_24_972 ();
 sg13g2_decap_8 FILLER_24_979 ();
 sg13g2_decap_8 FILLER_24_986 ();
 sg13g2_decap_8 FILLER_24_993 ();
 sg13g2_decap_8 FILLER_24_1000 ();
 sg13g2_decap_8 FILLER_24_1007 ();
 sg13g2_decap_8 FILLER_24_1014 ();
 sg13g2_decap_8 FILLER_24_1021 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_4 FILLER_25_32 ();
 sg13g2_fill_1 FILLER_25_63 ();
 sg13g2_fill_2 FILLER_25_69 ();
 sg13g2_fill_1 FILLER_25_71 ();
 sg13g2_decap_4 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_135 ();
 sg13g2_decap_4 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_146 ();
 sg13g2_decap_8 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_227 ();
 sg13g2_fill_2 FILLER_25_242 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_fill_2 FILLER_25_318 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_329 ();
 sg13g2_decap_4 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_4 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_424 ();
 sg13g2_decap_8 FILLER_25_431 ();
 sg13g2_fill_1 FILLER_25_438 ();
 sg13g2_decap_8 FILLER_25_443 ();
 sg13g2_decap_8 FILLER_25_450 ();
 sg13g2_decap_8 FILLER_25_457 ();
 sg13g2_decap_8 FILLER_25_464 ();
 sg13g2_decap_8 FILLER_25_471 ();
 sg13g2_decap_8 FILLER_25_478 ();
 sg13g2_decap_8 FILLER_25_485 ();
 sg13g2_decap_8 FILLER_25_492 ();
 sg13g2_decap_8 FILLER_25_499 ();
 sg13g2_decap_8 FILLER_25_506 ();
 sg13g2_decap_8 FILLER_25_513 ();
 sg13g2_decap_8 FILLER_25_520 ();
 sg13g2_decap_8 FILLER_25_527 ();
 sg13g2_decap_8 FILLER_25_534 ();
 sg13g2_decap_8 FILLER_25_541 ();
 sg13g2_decap_8 FILLER_25_548 ();
 sg13g2_decap_8 FILLER_25_555 ();
 sg13g2_decap_8 FILLER_25_562 ();
 sg13g2_decap_8 FILLER_25_569 ();
 sg13g2_decap_8 FILLER_25_576 ();
 sg13g2_decap_8 FILLER_25_583 ();
 sg13g2_decap_8 FILLER_25_590 ();
 sg13g2_decap_8 FILLER_25_597 ();
 sg13g2_decap_8 FILLER_25_604 ();
 sg13g2_decap_8 FILLER_25_611 ();
 sg13g2_decap_8 FILLER_25_618 ();
 sg13g2_decap_8 FILLER_25_625 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_decap_8 FILLER_25_639 ();
 sg13g2_decap_8 FILLER_25_646 ();
 sg13g2_decap_8 FILLER_25_653 ();
 sg13g2_decap_8 FILLER_25_660 ();
 sg13g2_decap_8 FILLER_25_667 ();
 sg13g2_decap_8 FILLER_25_674 ();
 sg13g2_decap_8 FILLER_25_681 ();
 sg13g2_decap_8 FILLER_25_688 ();
 sg13g2_decap_8 FILLER_25_695 ();
 sg13g2_decap_8 FILLER_25_702 ();
 sg13g2_decap_8 FILLER_25_709 ();
 sg13g2_decap_8 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_decap_8 FILLER_25_730 ();
 sg13g2_decap_8 FILLER_25_737 ();
 sg13g2_decap_8 FILLER_25_744 ();
 sg13g2_decap_8 FILLER_25_751 ();
 sg13g2_decap_8 FILLER_25_758 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_8 FILLER_25_856 ();
 sg13g2_decap_8 FILLER_25_863 ();
 sg13g2_decap_8 FILLER_25_870 ();
 sg13g2_decap_8 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_25_884 ();
 sg13g2_decap_8 FILLER_25_891 ();
 sg13g2_decap_8 FILLER_25_898 ();
 sg13g2_decap_8 FILLER_25_905 ();
 sg13g2_decap_8 FILLER_25_912 ();
 sg13g2_decap_8 FILLER_25_919 ();
 sg13g2_decap_8 FILLER_25_926 ();
 sg13g2_decap_8 FILLER_25_933 ();
 sg13g2_decap_8 FILLER_25_940 ();
 sg13g2_decap_8 FILLER_25_947 ();
 sg13g2_decap_8 FILLER_25_954 ();
 sg13g2_decap_8 FILLER_25_961 ();
 sg13g2_decap_8 FILLER_25_968 ();
 sg13g2_decap_8 FILLER_25_975 ();
 sg13g2_decap_8 FILLER_25_982 ();
 sg13g2_decap_8 FILLER_25_989 ();
 sg13g2_decap_8 FILLER_25_996 ();
 sg13g2_decap_8 FILLER_25_1003 ();
 sg13g2_decap_8 FILLER_25_1010 ();
 sg13g2_decap_8 FILLER_25_1017 ();
 sg13g2_decap_4 FILLER_25_1024 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_fill_2 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_82 ();
 sg13g2_fill_1 FILLER_26_92 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_decap_4 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_129 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_165 ();
 sg13g2_decap_4 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_4 FILLER_26_335 ();
 sg13g2_decap_4 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_4 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_fill_2 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_26_461 ();
 sg13g2_decap_8 FILLER_26_468 ();
 sg13g2_decap_8 FILLER_26_475 ();
 sg13g2_decap_8 FILLER_26_482 ();
 sg13g2_decap_8 FILLER_26_489 ();
 sg13g2_decap_8 FILLER_26_496 ();
 sg13g2_decap_8 FILLER_26_503 ();
 sg13g2_decap_8 FILLER_26_510 ();
 sg13g2_decap_8 FILLER_26_517 ();
 sg13g2_decap_8 FILLER_26_524 ();
 sg13g2_decap_8 FILLER_26_531 ();
 sg13g2_decap_8 FILLER_26_538 ();
 sg13g2_decap_8 FILLER_26_545 ();
 sg13g2_decap_8 FILLER_26_552 ();
 sg13g2_decap_8 FILLER_26_559 ();
 sg13g2_decap_8 FILLER_26_566 ();
 sg13g2_decap_8 FILLER_26_573 ();
 sg13g2_decap_8 FILLER_26_580 ();
 sg13g2_decap_8 FILLER_26_587 ();
 sg13g2_decap_8 FILLER_26_594 ();
 sg13g2_decap_8 FILLER_26_601 ();
 sg13g2_decap_8 FILLER_26_608 ();
 sg13g2_decap_8 FILLER_26_615 ();
 sg13g2_decap_8 FILLER_26_622 ();
 sg13g2_decap_8 FILLER_26_629 ();
 sg13g2_decap_8 FILLER_26_636 ();
 sg13g2_decap_8 FILLER_26_643 ();
 sg13g2_decap_8 FILLER_26_650 ();
 sg13g2_decap_8 FILLER_26_657 ();
 sg13g2_decap_8 FILLER_26_664 ();
 sg13g2_decap_8 FILLER_26_671 ();
 sg13g2_decap_8 FILLER_26_678 ();
 sg13g2_decap_8 FILLER_26_685 ();
 sg13g2_decap_8 FILLER_26_692 ();
 sg13g2_decap_8 FILLER_26_699 ();
 sg13g2_decap_8 FILLER_26_706 ();
 sg13g2_decap_8 FILLER_26_713 ();
 sg13g2_decap_8 FILLER_26_720 ();
 sg13g2_decap_8 FILLER_26_727 ();
 sg13g2_decap_8 FILLER_26_734 ();
 sg13g2_decap_8 FILLER_26_741 ();
 sg13g2_decap_8 FILLER_26_748 ();
 sg13g2_decap_8 FILLER_26_755 ();
 sg13g2_decap_8 FILLER_26_762 ();
 sg13g2_decap_8 FILLER_26_769 ();
 sg13g2_decap_8 FILLER_26_776 ();
 sg13g2_decap_8 FILLER_26_783 ();
 sg13g2_decap_8 FILLER_26_790 ();
 sg13g2_decap_8 FILLER_26_797 ();
 sg13g2_decap_8 FILLER_26_804 ();
 sg13g2_decap_8 FILLER_26_811 ();
 sg13g2_decap_8 FILLER_26_818 ();
 sg13g2_decap_8 FILLER_26_825 ();
 sg13g2_decap_8 FILLER_26_832 ();
 sg13g2_decap_8 FILLER_26_839 ();
 sg13g2_decap_8 FILLER_26_846 ();
 sg13g2_decap_8 FILLER_26_853 ();
 sg13g2_decap_8 FILLER_26_860 ();
 sg13g2_decap_8 FILLER_26_867 ();
 sg13g2_decap_8 FILLER_26_874 ();
 sg13g2_decap_8 FILLER_26_881 ();
 sg13g2_decap_8 FILLER_26_888 ();
 sg13g2_decap_8 FILLER_26_895 ();
 sg13g2_decap_8 FILLER_26_902 ();
 sg13g2_decap_8 FILLER_26_909 ();
 sg13g2_decap_8 FILLER_26_916 ();
 sg13g2_decap_8 FILLER_26_923 ();
 sg13g2_decap_8 FILLER_26_930 ();
 sg13g2_decap_8 FILLER_26_937 ();
 sg13g2_decap_8 FILLER_26_944 ();
 sg13g2_decap_8 FILLER_26_951 ();
 sg13g2_decap_8 FILLER_26_958 ();
 sg13g2_decap_8 FILLER_26_965 ();
 sg13g2_decap_8 FILLER_26_972 ();
 sg13g2_decap_8 FILLER_26_979 ();
 sg13g2_decap_8 FILLER_26_986 ();
 sg13g2_decap_8 FILLER_26_993 ();
 sg13g2_decap_8 FILLER_26_1000 ();
 sg13g2_decap_8 FILLER_26_1007 ();
 sg13g2_decap_8 FILLER_26_1014 ();
 sg13g2_decap_8 FILLER_26_1021 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_15 ();
 sg13g2_fill_1 FILLER_27_20 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_decap_8 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_decap_4 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_405 ();
 sg13g2_fill_2 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_decap_8 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_decap_8 FILLER_27_889 ();
 sg13g2_decap_8 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_910 ();
 sg13g2_decap_8 FILLER_27_917 ();
 sg13g2_decap_8 FILLER_27_924 ();
 sg13g2_decap_8 FILLER_27_931 ();
 sg13g2_decap_8 FILLER_27_938 ();
 sg13g2_decap_8 FILLER_27_945 ();
 sg13g2_decap_8 FILLER_27_952 ();
 sg13g2_decap_8 FILLER_27_959 ();
 sg13g2_decap_8 FILLER_27_966 ();
 sg13g2_decap_8 FILLER_27_973 ();
 sg13g2_decap_8 FILLER_27_980 ();
 sg13g2_decap_8 FILLER_27_987 ();
 sg13g2_decap_8 FILLER_27_994 ();
 sg13g2_decap_8 FILLER_27_1001 ();
 sg13g2_decap_8 FILLER_27_1008 ();
 sg13g2_decap_8 FILLER_27_1015 ();
 sg13g2_decap_8 FILLER_27_1022 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_decap_4 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_117 ();
 sg13g2_fill_2 FILLER_28_132 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_170 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_decap_8 FILLER_28_223 ();
 sg13g2_decap_4 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_393 ();
 sg13g2_fill_1 FILLER_28_462 ();
 sg13g2_decap_4 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_508 ();
 sg13g2_decap_8 FILLER_28_515 ();
 sg13g2_decap_8 FILLER_28_522 ();
 sg13g2_decap_8 FILLER_28_529 ();
 sg13g2_decap_8 FILLER_28_536 ();
 sg13g2_decap_8 FILLER_28_543 ();
 sg13g2_decap_8 FILLER_28_550 ();
 sg13g2_decap_8 FILLER_28_557 ();
 sg13g2_decap_8 FILLER_28_564 ();
 sg13g2_decap_8 FILLER_28_571 ();
 sg13g2_decap_8 FILLER_28_578 ();
 sg13g2_decap_8 FILLER_28_585 ();
 sg13g2_decap_8 FILLER_28_592 ();
 sg13g2_decap_8 FILLER_28_599 ();
 sg13g2_decap_8 FILLER_28_606 ();
 sg13g2_decap_8 FILLER_28_613 ();
 sg13g2_decap_8 FILLER_28_620 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_decap_8 FILLER_28_634 ();
 sg13g2_decap_8 FILLER_28_641 ();
 sg13g2_decap_8 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_655 ();
 sg13g2_decap_8 FILLER_28_662 ();
 sg13g2_decap_8 FILLER_28_669 ();
 sg13g2_decap_8 FILLER_28_676 ();
 sg13g2_decap_8 FILLER_28_683 ();
 sg13g2_decap_8 FILLER_28_690 ();
 sg13g2_decap_8 FILLER_28_697 ();
 sg13g2_decap_8 FILLER_28_704 ();
 sg13g2_decap_8 FILLER_28_711 ();
 sg13g2_decap_8 FILLER_28_718 ();
 sg13g2_decap_8 FILLER_28_725 ();
 sg13g2_decap_8 FILLER_28_732 ();
 sg13g2_decap_8 FILLER_28_739 ();
 sg13g2_decap_8 FILLER_28_746 ();
 sg13g2_decap_8 FILLER_28_753 ();
 sg13g2_decap_8 FILLER_28_760 ();
 sg13g2_decap_8 FILLER_28_767 ();
 sg13g2_decap_8 FILLER_28_774 ();
 sg13g2_decap_8 FILLER_28_781 ();
 sg13g2_decap_8 FILLER_28_788 ();
 sg13g2_decap_8 FILLER_28_795 ();
 sg13g2_decap_8 FILLER_28_802 ();
 sg13g2_decap_8 FILLER_28_809 ();
 sg13g2_decap_8 FILLER_28_816 ();
 sg13g2_decap_8 FILLER_28_823 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_decap_8 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_28_865 ();
 sg13g2_decap_8 FILLER_28_872 ();
 sg13g2_decap_8 FILLER_28_879 ();
 sg13g2_decap_8 FILLER_28_886 ();
 sg13g2_decap_8 FILLER_28_893 ();
 sg13g2_decap_8 FILLER_28_900 ();
 sg13g2_decap_8 FILLER_28_907 ();
 sg13g2_decap_8 FILLER_28_914 ();
 sg13g2_decap_8 FILLER_28_921 ();
 sg13g2_decap_8 FILLER_28_928 ();
 sg13g2_decap_8 FILLER_28_935 ();
 sg13g2_decap_8 FILLER_28_942 ();
 sg13g2_decap_8 FILLER_28_949 ();
 sg13g2_decap_8 FILLER_28_956 ();
 sg13g2_decap_8 FILLER_28_963 ();
 sg13g2_decap_8 FILLER_28_970 ();
 sg13g2_decap_8 FILLER_28_977 ();
 sg13g2_decap_8 FILLER_28_984 ();
 sg13g2_decap_8 FILLER_28_991 ();
 sg13g2_decap_8 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1005 ();
 sg13g2_decap_8 FILLER_28_1012 ();
 sg13g2_decap_8 FILLER_28_1019 ();
 sg13g2_fill_2 FILLER_28_1026 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_fill_2 FILLER_29_4 ();
 sg13g2_fill_1 FILLER_29_33 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_59 ();
 sg13g2_decap_4 FILLER_29_85 ();
 sg13g2_decap_4 FILLER_29_103 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_decap_4 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_378 ();
 sg13g2_fill_1 FILLER_29_402 ();
 sg13g2_fill_2 FILLER_29_451 ();
 sg13g2_decap_8 FILLER_29_493 ();
 sg13g2_decap_8 FILLER_29_528 ();
 sg13g2_decap_8 FILLER_29_535 ();
 sg13g2_decap_8 FILLER_29_542 ();
 sg13g2_decap_8 FILLER_29_549 ();
 sg13g2_decap_8 FILLER_29_556 ();
 sg13g2_decap_8 FILLER_29_563 ();
 sg13g2_decap_8 FILLER_29_570 ();
 sg13g2_decap_8 FILLER_29_577 ();
 sg13g2_decap_8 FILLER_29_584 ();
 sg13g2_decap_8 FILLER_29_591 ();
 sg13g2_decap_8 FILLER_29_598 ();
 sg13g2_decap_8 FILLER_29_605 ();
 sg13g2_decap_8 FILLER_29_612 ();
 sg13g2_decap_8 FILLER_29_619 ();
 sg13g2_decap_8 FILLER_29_626 ();
 sg13g2_decap_8 FILLER_29_633 ();
 sg13g2_decap_8 FILLER_29_640 ();
 sg13g2_decap_8 FILLER_29_647 ();
 sg13g2_decap_8 FILLER_29_654 ();
 sg13g2_decap_8 FILLER_29_661 ();
 sg13g2_decap_8 FILLER_29_668 ();
 sg13g2_decap_8 FILLER_29_675 ();
 sg13g2_decap_8 FILLER_29_682 ();
 sg13g2_decap_8 FILLER_29_689 ();
 sg13g2_decap_8 FILLER_29_696 ();
 sg13g2_decap_8 FILLER_29_703 ();
 sg13g2_decap_8 FILLER_29_710 ();
 sg13g2_decap_8 FILLER_29_717 ();
 sg13g2_decap_8 FILLER_29_724 ();
 sg13g2_decap_8 FILLER_29_731 ();
 sg13g2_decap_8 FILLER_29_738 ();
 sg13g2_decap_8 FILLER_29_745 ();
 sg13g2_decap_8 FILLER_29_752 ();
 sg13g2_decap_8 FILLER_29_759 ();
 sg13g2_decap_8 FILLER_29_766 ();
 sg13g2_decap_8 FILLER_29_773 ();
 sg13g2_decap_8 FILLER_29_780 ();
 sg13g2_decap_8 FILLER_29_787 ();
 sg13g2_decap_8 FILLER_29_794 ();
 sg13g2_decap_8 FILLER_29_801 ();
 sg13g2_decap_8 FILLER_29_808 ();
 sg13g2_decap_8 FILLER_29_815 ();
 sg13g2_decap_8 FILLER_29_822 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_decap_8 FILLER_29_836 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_850 ();
 sg13g2_decap_8 FILLER_29_857 ();
 sg13g2_decap_8 FILLER_29_864 ();
 sg13g2_decap_8 FILLER_29_871 ();
 sg13g2_decap_8 FILLER_29_878 ();
 sg13g2_decap_8 FILLER_29_885 ();
 sg13g2_decap_8 FILLER_29_892 ();
 sg13g2_decap_8 FILLER_29_899 ();
 sg13g2_decap_8 FILLER_29_906 ();
 sg13g2_decap_8 FILLER_29_913 ();
 sg13g2_decap_8 FILLER_29_920 ();
 sg13g2_decap_8 FILLER_29_927 ();
 sg13g2_decap_8 FILLER_29_934 ();
 sg13g2_decap_8 FILLER_29_941 ();
 sg13g2_decap_8 FILLER_29_948 ();
 sg13g2_decap_8 FILLER_29_955 ();
 sg13g2_decap_8 FILLER_29_962 ();
 sg13g2_decap_8 FILLER_29_969 ();
 sg13g2_decap_8 FILLER_29_976 ();
 sg13g2_decap_8 FILLER_29_983 ();
 sg13g2_decap_8 FILLER_29_990 ();
 sg13g2_decap_8 FILLER_29_997 ();
 sg13g2_decap_8 FILLER_29_1004 ();
 sg13g2_decap_8 FILLER_29_1011 ();
 sg13g2_decap_8 FILLER_29_1018 ();
 sg13g2_decap_4 FILLER_29_1025 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_15 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_decap_8 FILLER_30_184 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_decap_4 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_decap_4 FILLER_30_322 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_fill_1 FILLER_30_420 ();
 sg13g2_fill_2 FILLER_30_486 ();
 sg13g2_fill_1 FILLER_30_488 ();
 sg13g2_fill_2 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_517 ();
 sg13g2_decap_8 FILLER_30_524 ();
 sg13g2_decap_8 FILLER_30_531 ();
 sg13g2_decap_8 FILLER_30_538 ();
 sg13g2_decap_8 FILLER_30_545 ();
 sg13g2_decap_8 FILLER_30_552 ();
 sg13g2_decap_8 FILLER_30_559 ();
 sg13g2_decap_8 FILLER_30_566 ();
 sg13g2_decap_8 FILLER_30_573 ();
 sg13g2_decap_8 FILLER_30_580 ();
 sg13g2_decap_8 FILLER_30_587 ();
 sg13g2_decap_8 FILLER_30_594 ();
 sg13g2_decap_8 FILLER_30_601 ();
 sg13g2_decap_8 FILLER_30_608 ();
 sg13g2_decap_8 FILLER_30_615 ();
 sg13g2_decap_8 FILLER_30_622 ();
 sg13g2_decap_8 FILLER_30_629 ();
 sg13g2_decap_8 FILLER_30_636 ();
 sg13g2_decap_8 FILLER_30_643 ();
 sg13g2_decap_8 FILLER_30_650 ();
 sg13g2_decap_8 FILLER_30_657 ();
 sg13g2_decap_8 FILLER_30_664 ();
 sg13g2_decap_8 FILLER_30_671 ();
 sg13g2_decap_8 FILLER_30_678 ();
 sg13g2_decap_8 FILLER_30_685 ();
 sg13g2_decap_8 FILLER_30_692 ();
 sg13g2_decap_8 FILLER_30_699 ();
 sg13g2_decap_8 FILLER_30_706 ();
 sg13g2_decap_8 FILLER_30_713 ();
 sg13g2_decap_8 FILLER_30_720 ();
 sg13g2_decap_8 FILLER_30_727 ();
 sg13g2_decap_8 FILLER_30_734 ();
 sg13g2_decap_8 FILLER_30_741 ();
 sg13g2_decap_8 FILLER_30_748 ();
 sg13g2_decap_8 FILLER_30_755 ();
 sg13g2_decap_8 FILLER_30_762 ();
 sg13g2_decap_8 FILLER_30_769 ();
 sg13g2_decap_8 FILLER_30_776 ();
 sg13g2_decap_8 FILLER_30_783 ();
 sg13g2_decap_8 FILLER_30_790 ();
 sg13g2_decap_8 FILLER_30_797 ();
 sg13g2_decap_8 FILLER_30_804 ();
 sg13g2_decap_8 FILLER_30_811 ();
 sg13g2_decap_8 FILLER_30_818 ();
 sg13g2_decap_8 FILLER_30_825 ();
 sg13g2_decap_8 FILLER_30_832 ();
 sg13g2_decap_8 FILLER_30_839 ();
 sg13g2_decap_8 FILLER_30_846 ();
 sg13g2_decap_8 FILLER_30_853 ();
 sg13g2_decap_8 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_30_867 ();
 sg13g2_decap_8 FILLER_30_874 ();
 sg13g2_decap_8 FILLER_30_881 ();
 sg13g2_decap_8 FILLER_30_888 ();
 sg13g2_decap_8 FILLER_30_895 ();
 sg13g2_decap_8 FILLER_30_902 ();
 sg13g2_decap_8 FILLER_30_909 ();
 sg13g2_decap_8 FILLER_30_916 ();
 sg13g2_decap_8 FILLER_30_923 ();
 sg13g2_decap_8 FILLER_30_930 ();
 sg13g2_decap_8 FILLER_30_937 ();
 sg13g2_decap_8 FILLER_30_944 ();
 sg13g2_decap_8 FILLER_30_951 ();
 sg13g2_decap_8 FILLER_30_958 ();
 sg13g2_decap_8 FILLER_30_965 ();
 sg13g2_decap_8 FILLER_30_972 ();
 sg13g2_decap_8 FILLER_30_979 ();
 sg13g2_decap_8 FILLER_30_986 ();
 sg13g2_decap_8 FILLER_30_993 ();
 sg13g2_decap_8 FILLER_30_1000 ();
 sg13g2_decap_8 FILLER_30_1007 ();
 sg13g2_decap_8 FILLER_30_1014 ();
 sg13g2_decap_8 FILLER_30_1021 ();
 sg13g2_fill_1 FILLER_30_1028 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_decap_4 FILLER_31_32 ();
 sg13g2_decap_4 FILLER_31_92 ();
 sg13g2_fill_2 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_decap_4 FILLER_31_182 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_247 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_279 ();
 sg13g2_decap_4 FILLER_31_293 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_31_326 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_372 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_2 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_402 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_2 FILLER_31_429 ();
 sg13g2_fill_1 FILLER_31_431 ();
 sg13g2_fill_1 FILLER_31_449 ();
 sg13g2_fill_1 FILLER_31_492 ();
 sg13g2_fill_2 FILLER_31_506 ();
 sg13g2_decap_8 FILLER_31_536 ();
 sg13g2_decap_8 FILLER_31_543 ();
 sg13g2_decap_8 FILLER_31_550 ();
 sg13g2_decap_8 FILLER_31_557 ();
 sg13g2_decap_8 FILLER_31_564 ();
 sg13g2_decap_8 FILLER_31_571 ();
 sg13g2_decap_8 FILLER_31_578 ();
 sg13g2_decap_8 FILLER_31_585 ();
 sg13g2_decap_8 FILLER_31_592 ();
 sg13g2_decap_8 FILLER_31_599 ();
 sg13g2_decap_8 FILLER_31_606 ();
 sg13g2_decap_8 FILLER_31_613 ();
 sg13g2_decap_8 FILLER_31_620 ();
 sg13g2_decap_8 FILLER_31_627 ();
 sg13g2_decap_8 FILLER_31_634 ();
 sg13g2_decap_8 FILLER_31_641 ();
 sg13g2_decap_8 FILLER_31_648 ();
 sg13g2_decap_8 FILLER_31_655 ();
 sg13g2_decap_8 FILLER_31_662 ();
 sg13g2_decap_8 FILLER_31_669 ();
 sg13g2_decap_8 FILLER_31_676 ();
 sg13g2_decap_8 FILLER_31_683 ();
 sg13g2_decap_8 FILLER_31_690 ();
 sg13g2_decap_8 FILLER_31_697 ();
 sg13g2_decap_8 FILLER_31_704 ();
 sg13g2_decap_8 FILLER_31_711 ();
 sg13g2_decap_8 FILLER_31_718 ();
 sg13g2_decap_8 FILLER_31_725 ();
 sg13g2_decap_8 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_739 ();
 sg13g2_decap_8 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_753 ();
 sg13g2_decap_8 FILLER_31_760 ();
 sg13g2_decap_8 FILLER_31_767 ();
 sg13g2_decap_8 FILLER_31_774 ();
 sg13g2_decap_8 FILLER_31_781 ();
 sg13g2_decap_8 FILLER_31_788 ();
 sg13g2_decap_8 FILLER_31_795 ();
 sg13g2_decap_8 FILLER_31_802 ();
 sg13g2_decap_8 FILLER_31_809 ();
 sg13g2_decap_8 FILLER_31_816 ();
 sg13g2_decap_8 FILLER_31_823 ();
 sg13g2_decap_8 FILLER_31_830 ();
 sg13g2_decap_8 FILLER_31_837 ();
 sg13g2_decap_8 FILLER_31_844 ();
 sg13g2_decap_8 FILLER_31_851 ();
 sg13g2_decap_8 FILLER_31_858 ();
 sg13g2_decap_8 FILLER_31_865 ();
 sg13g2_decap_8 FILLER_31_872 ();
 sg13g2_decap_8 FILLER_31_879 ();
 sg13g2_decap_8 FILLER_31_886 ();
 sg13g2_decap_8 FILLER_31_893 ();
 sg13g2_decap_8 FILLER_31_900 ();
 sg13g2_decap_8 FILLER_31_907 ();
 sg13g2_decap_8 FILLER_31_914 ();
 sg13g2_decap_8 FILLER_31_921 ();
 sg13g2_decap_8 FILLER_31_928 ();
 sg13g2_decap_8 FILLER_31_935 ();
 sg13g2_decap_8 FILLER_31_942 ();
 sg13g2_decap_8 FILLER_31_949 ();
 sg13g2_decap_8 FILLER_31_956 ();
 sg13g2_decap_8 FILLER_31_963 ();
 sg13g2_decap_8 FILLER_31_970 ();
 sg13g2_decap_8 FILLER_31_977 ();
 sg13g2_decap_8 FILLER_31_984 ();
 sg13g2_decap_8 FILLER_31_991 ();
 sg13g2_decap_8 FILLER_31_998 ();
 sg13g2_decap_8 FILLER_31_1005 ();
 sg13g2_decap_8 FILLER_31_1012 ();
 sg13g2_decap_8 FILLER_31_1019 ();
 sg13g2_fill_2 FILLER_31_1026 ();
 sg13g2_fill_1 FILLER_31_1028 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_69 ();
 sg13g2_fill_2 FILLER_32_73 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_303 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_315 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_fill_1 FILLER_32_398 ();
 sg13g2_fill_2 FILLER_32_420 ();
 sg13g2_fill_1 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_433 ();
 sg13g2_fill_2 FILLER_32_447 ();
 sg13g2_fill_1 FILLER_32_454 ();
 sg13g2_decap_8 FILLER_32_528 ();
 sg13g2_decap_8 FILLER_32_535 ();
 sg13g2_decap_8 FILLER_32_542 ();
 sg13g2_decap_8 FILLER_32_549 ();
 sg13g2_decap_8 FILLER_32_556 ();
 sg13g2_decap_8 FILLER_32_563 ();
 sg13g2_decap_8 FILLER_32_570 ();
 sg13g2_decap_8 FILLER_32_577 ();
 sg13g2_decap_8 FILLER_32_584 ();
 sg13g2_decap_8 FILLER_32_591 ();
 sg13g2_decap_8 FILLER_32_598 ();
 sg13g2_decap_8 FILLER_32_605 ();
 sg13g2_decap_8 FILLER_32_612 ();
 sg13g2_decap_8 FILLER_32_619 ();
 sg13g2_decap_8 FILLER_32_626 ();
 sg13g2_decap_8 FILLER_32_633 ();
 sg13g2_decap_8 FILLER_32_640 ();
 sg13g2_decap_8 FILLER_32_647 ();
 sg13g2_decap_8 FILLER_32_654 ();
 sg13g2_decap_8 FILLER_32_661 ();
 sg13g2_decap_8 FILLER_32_668 ();
 sg13g2_decap_8 FILLER_32_675 ();
 sg13g2_decap_8 FILLER_32_682 ();
 sg13g2_decap_8 FILLER_32_689 ();
 sg13g2_decap_8 FILLER_32_696 ();
 sg13g2_decap_8 FILLER_32_703 ();
 sg13g2_decap_8 FILLER_32_710 ();
 sg13g2_decap_8 FILLER_32_717 ();
 sg13g2_decap_8 FILLER_32_724 ();
 sg13g2_decap_8 FILLER_32_731 ();
 sg13g2_decap_8 FILLER_32_738 ();
 sg13g2_decap_8 FILLER_32_745 ();
 sg13g2_decap_8 FILLER_32_752 ();
 sg13g2_decap_8 FILLER_32_759 ();
 sg13g2_decap_8 FILLER_32_766 ();
 sg13g2_decap_8 FILLER_32_773 ();
 sg13g2_decap_8 FILLER_32_780 ();
 sg13g2_decap_8 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_794 ();
 sg13g2_decap_8 FILLER_32_801 ();
 sg13g2_decap_8 FILLER_32_808 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_decap_8 FILLER_32_822 ();
 sg13g2_decap_8 FILLER_32_829 ();
 sg13g2_decap_8 FILLER_32_836 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_decap_8 FILLER_32_864 ();
 sg13g2_decap_8 FILLER_32_871 ();
 sg13g2_decap_8 FILLER_32_878 ();
 sg13g2_decap_8 FILLER_32_885 ();
 sg13g2_decap_8 FILLER_32_892 ();
 sg13g2_decap_8 FILLER_32_899 ();
 sg13g2_decap_8 FILLER_32_906 ();
 sg13g2_decap_8 FILLER_32_913 ();
 sg13g2_decap_8 FILLER_32_920 ();
 sg13g2_decap_8 FILLER_32_927 ();
 sg13g2_decap_8 FILLER_32_934 ();
 sg13g2_decap_8 FILLER_32_941 ();
 sg13g2_decap_8 FILLER_32_948 ();
 sg13g2_decap_8 FILLER_32_955 ();
 sg13g2_decap_8 FILLER_32_962 ();
 sg13g2_decap_8 FILLER_32_969 ();
 sg13g2_decap_8 FILLER_32_976 ();
 sg13g2_decap_8 FILLER_32_983 ();
 sg13g2_decap_8 FILLER_32_990 ();
 sg13g2_decap_8 FILLER_32_997 ();
 sg13g2_decap_8 FILLER_32_1004 ();
 sg13g2_decap_8 FILLER_32_1011 ();
 sg13g2_decap_8 FILLER_32_1018 ();
 sg13g2_decap_4 FILLER_32_1025 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_43 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_decap_4 FILLER_33_80 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_fill_2 FILLER_33_179 ();
 sg13g2_fill_1 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_decap_4 FILLER_33_284 ();
 sg13g2_decap_4 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_332 ();
 sg13g2_decap_4 FILLER_33_339 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_decap_4 FILLER_33_395 ();
 sg13g2_fill_2 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_decap_4 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_33_438 ();
 sg13g2_fill_2 FILLER_33_452 ();
 sg13g2_fill_2 FILLER_33_463 ();
 sg13g2_fill_2 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_533 ();
 sg13g2_decap_8 FILLER_33_540 ();
 sg13g2_decap_8 FILLER_33_547 ();
 sg13g2_decap_8 FILLER_33_554 ();
 sg13g2_decap_8 FILLER_33_561 ();
 sg13g2_decap_8 FILLER_33_568 ();
 sg13g2_decap_8 FILLER_33_575 ();
 sg13g2_decap_8 FILLER_33_582 ();
 sg13g2_decap_8 FILLER_33_589 ();
 sg13g2_decap_8 FILLER_33_596 ();
 sg13g2_decap_8 FILLER_33_603 ();
 sg13g2_decap_8 FILLER_33_610 ();
 sg13g2_decap_8 FILLER_33_617 ();
 sg13g2_decap_8 FILLER_33_624 ();
 sg13g2_decap_8 FILLER_33_631 ();
 sg13g2_decap_8 FILLER_33_638 ();
 sg13g2_decap_8 FILLER_33_645 ();
 sg13g2_decap_8 FILLER_33_652 ();
 sg13g2_decap_8 FILLER_33_659 ();
 sg13g2_decap_8 FILLER_33_666 ();
 sg13g2_decap_8 FILLER_33_673 ();
 sg13g2_decap_8 FILLER_33_680 ();
 sg13g2_decap_8 FILLER_33_687 ();
 sg13g2_decap_8 FILLER_33_694 ();
 sg13g2_decap_8 FILLER_33_701 ();
 sg13g2_decap_8 FILLER_33_708 ();
 sg13g2_decap_8 FILLER_33_715 ();
 sg13g2_decap_8 FILLER_33_722 ();
 sg13g2_decap_8 FILLER_33_729 ();
 sg13g2_decap_8 FILLER_33_736 ();
 sg13g2_decap_8 FILLER_33_743 ();
 sg13g2_decap_8 FILLER_33_750 ();
 sg13g2_decap_8 FILLER_33_757 ();
 sg13g2_decap_8 FILLER_33_764 ();
 sg13g2_decap_8 FILLER_33_771 ();
 sg13g2_decap_8 FILLER_33_778 ();
 sg13g2_decap_8 FILLER_33_785 ();
 sg13g2_decap_8 FILLER_33_792 ();
 sg13g2_decap_8 FILLER_33_799 ();
 sg13g2_decap_8 FILLER_33_806 ();
 sg13g2_decap_8 FILLER_33_813 ();
 sg13g2_decap_8 FILLER_33_820 ();
 sg13g2_decap_8 FILLER_33_827 ();
 sg13g2_decap_8 FILLER_33_834 ();
 sg13g2_decap_8 FILLER_33_841 ();
 sg13g2_decap_8 FILLER_33_848 ();
 sg13g2_decap_8 FILLER_33_855 ();
 sg13g2_decap_8 FILLER_33_862 ();
 sg13g2_decap_8 FILLER_33_869 ();
 sg13g2_decap_8 FILLER_33_876 ();
 sg13g2_decap_8 FILLER_33_883 ();
 sg13g2_decap_8 FILLER_33_890 ();
 sg13g2_decap_8 FILLER_33_897 ();
 sg13g2_decap_8 FILLER_33_904 ();
 sg13g2_decap_8 FILLER_33_911 ();
 sg13g2_decap_8 FILLER_33_918 ();
 sg13g2_decap_8 FILLER_33_925 ();
 sg13g2_decap_8 FILLER_33_932 ();
 sg13g2_decap_8 FILLER_33_939 ();
 sg13g2_decap_8 FILLER_33_946 ();
 sg13g2_decap_8 FILLER_33_953 ();
 sg13g2_decap_8 FILLER_33_960 ();
 sg13g2_decap_8 FILLER_33_967 ();
 sg13g2_decap_8 FILLER_33_974 ();
 sg13g2_decap_8 FILLER_33_981 ();
 sg13g2_decap_8 FILLER_33_988 ();
 sg13g2_decap_8 FILLER_33_995 ();
 sg13g2_decap_8 FILLER_33_1002 ();
 sg13g2_decap_8 FILLER_33_1009 ();
 sg13g2_decap_8 FILLER_33_1016 ();
 sg13g2_decap_4 FILLER_33_1023 ();
 sg13g2_fill_2 FILLER_33_1027 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_69 ();
 sg13g2_fill_1 FILLER_34_71 ();
 sg13g2_decap_4 FILLER_34_85 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_decap_4 FILLER_34_162 ();
 sg13g2_fill_2 FILLER_34_166 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_decap_8 FILLER_34_235 ();
 sg13g2_decap_4 FILLER_34_242 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_decap_4 FILLER_34_270 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_decap_4 FILLER_34_289 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_304 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_408 ();
 sg13g2_fill_1 FILLER_34_410 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_decap_4 FILLER_34_464 ();
 sg13g2_fill_1 FILLER_34_509 ();
 sg13g2_decap_8 FILLER_34_537 ();
 sg13g2_decap_8 FILLER_34_544 ();
 sg13g2_decap_8 FILLER_34_551 ();
 sg13g2_decap_8 FILLER_34_558 ();
 sg13g2_decap_8 FILLER_34_565 ();
 sg13g2_decap_8 FILLER_34_572 ();
 sg13g2_decap_8 FILLER_34_579 ();
 sg13g2_decap_8 FILLER_34_586 ();
 sg13g2_decap_8 FILLER_34_593 ();
 sg13g2_decap_8 FILLER_34_600 ();
 sg13g2_decap_8 FILLER_34_607 ();
 sg13g2_decap_8 FILLER_34_614 ();
 sg13g2_decap_8 FILLER_34_621 ();
 sg13g2_decap_8 FILLER_34_628 ();
 sg13g2_decap_8 FILLER_34_635 ();
 sg13g2_decap_8 FILLER_34_642 ();
 sg13g2_decap_8 FILLER_34_649 ();
 sg13g2_decap_8 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_663 ();
 sg13g2_decap_8 FILLER_34_670 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_691 ();
 sg13g2_decap_8 FILLER_34_698 ();
 sg13g2_decap_8 FILLER_34_705 ();
 sg13g2_decap_8 FILLER_34_712 ();
 sg13g2_decap_8 FILLER_34_719 ();
 sg13g2_decap_8 FILLER_34_726 ();
 sg13g2_decap_8 FILLER_34_733 ();
 sg13g2_decap_8 FILLER_34_740 ();
 sg13g2_decap_8 FILLER_34_747 ();
 sg13g2_decap_8 FILLER_34_754 ();
 sg13g2_decap_8 FILLER_34_761 ();
 sg13g2_decap_8 FILLER_34_768 ();
 sg13g2_decap_8 FILLER_34_775 ();
 sg13g2_decap_8 FILLER_34_782 ();
 sg13g2_decap_8 FILLER_34_789 ();
 sg13g2_decap_8 FILLER_34_796 ();
 sg13g2_decap_8 FILLER_34_803 ();
 sg13g2_decap_8 FILLER_34_810 ();
 sg13g2_decap_8 FILLER_34_817 ();
 sg13g2_decap_8 FILLER_34_824 ();
 sg13g2_decap_8 FILLER_34_831 ();
 sg13g2_decap_8 FILLER_34_838 ();
 sg13g2_decap_8 FILLER_34_845 ();
 sg13g2_decap_8 FILLER_34_852 ();
 sg13g2_decap_8 FILLER_34_859 ();
 sg13g2_decap_8 FILLER_34_866 ();
 sg13g2_decap_8 FILLER_34_873 ();
 sg13g2_decap_8 FILLER_34_880 ();
 sg13g2_decap_8 FILLER_34_887 ();
 sg13g2_decap_8 FILLER_34_894 ();
 sg13g2_decap_8 FILLER_34_901 ();
 sg13g2_decap_8 FILLER_34_908 ();
 sg13g2_decap_8 FILLER_34_915 ();
 sg13g2_decap_8 FILLER_34_922 ();
 sg13g2_decap_8 FILLER_34_929 ();
 sg13g2_decap_8 FILLER_34_936 ();
 sg13g2_decap_8 FILLER_34_943 ();
 sg13g2_decap_8 FILLER_34_950 ();
 sg13g2_decap_8 FILLER_34_957 ();
 sg13g2_decap_8 FILLER_34_964 ();
 sg13g2_decap_8 FILLER_34_971 ();
 sg13g2_decap_8 FILLER_34_978 ();
 sg13g2_decap_8 FILLER_34_985 ();
 sg13g2_decap_8 FILLER_34_992 ();
 sg13g2_decap_8 FILLER_34_999 ();
 sg13g2_decap_8 FILLER_34_1006 ();
 sg13g2_decap_8 FILLER_34_1013 ();
 sg13g2_decap_8 FILLER_34_1020 ();
 sg13g2_fill_2 FILLER_34_1027 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_15 ();
 sg13g2_fill_2 FILLER_35_19 ();
 sg13g2_fill_1 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_128 ();
 sg13g2_decap_4 FILLER_35_143 ();
 sg13g2_decap_4 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_159 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_172 ();
 sg13g2_decap_4 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_decap_4 FILLER_35_305 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_decap_4 FILLER_35_330 ();
 sg13g2_fill_2 FILLER_35_334 ();
 sg13g2_decap_4 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_decap_4 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_396 ();
 sg13g2_fill_1 FILLER_35_398 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_414 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_decap_4 FILLER_35_428 ();
 sg13g2_fill_1 FILLER_35_432 ();
 sg13g2_fill_2 FILLER_35_437 ();
 sg13g2_fill_1 FILLER_35_439 ();
 sg13g2_fill_2 FILLER_35_453 ();
 sg13g2_decap_4 FILLER_35_459 ();
 sg13g2_decap_4 FILLER_35_468 ();
 sg13g2_fill_1 FILLER_35_481 ();
 sg13g2_fill_2 FILLER_35_493 ();
 sg13g2_fill_1 FILLER_35_505 ();
 sg13g2_decap_8 FILLER_35_533 ();
 sg13g2_decap_8 FILLER_35_540 ();
 sg13g2_decap_8 FILLER_35_547 ();
 sg13g2_decap_8 FILLER_35_554 ();
 sg13g2_decap_8 FILLER_35_561 ();
 sg13g2_decap_8 FILLER_35_568 ();
 sg13g2_decap_8 FILLER_35_575 ();
 sg13g2_decap_8 FILLER_35_582 ();
 sg13g2_decap_8 FILLER_35_589 ();
 sg13g2_decap_8 FILLER_35_596 ();
 sg13g2_decap_8 FILLER_35_603 ();
 sg13g2_decap_8 FILLER_35_610 ();
 sg13g2_decap_8 FILLER_35_617 ();
 sg13g2_decap_8 FILLER_35_624 ();
 sg13g2_decap_8 FILLER_35_631 ();
 sg13g2_decap_8 FILLER_35_638 ();
 sg13g2_decap_8 FILLER_35_645 ();
 sg13g2_decap_8 FILLER_35_652 ();
 sg13g2_decap_8 FILLER_35_659 ();
 sg13g2_decap_8 FILLER_35_666 ();
 sg13g2_decap_8 FILLER_35_673 ();
 sg13g2_decap_8 FILLER_35_680 ();
 sg13g2_decap_8 FILLER_35_687 ();
 sg13g2_decap_8 FILLER_35_694 ();
 sg13g2_decap_8 FILLER_35_701 ();
 sg13g2_decap_8 FILLER_35_708 ();
 sg13g2_decap_8 FILLER_35_715 ();
 sg13g2_decap_8 FILLER_35_722 ();
 sg13g2_decap_8 FILLER_35_729 ();
 sg13g2_decap_8 FILLER_35_736 ();
 sg13g2_decap_8 FILLER_35_743 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_decap_8 FILLER_35_757 ();
 sg13g2_decap_8 FILLER_35_764 ();
 sg13g2_decap_8 FILLER_35_771 ();
 sg13g2_decap_8 FILLER_35_778 ();
 sg13g2_decap_8 FILLER_35_785 ();
 sg13g2_decap_8 FILLER_35_792 ();
 sg13g2_decap_8 FILLER_35_799 ();
 sg13g2_decap_8 FILLER_35_806 ();
 sg13g2_decap_8 FILLER_35_813 ();
 sg13g2_decap_8 FILLER_35_820 ();
 sg13g2_decap_8 FILLER_35_827 ();
 sg13g2_decap_8 FILLER_35_834 ();
 sg13g2_decap_8 FILLER_35_841 ();
 sg13g2_decap_8 FILLER_35_848 ();
 sg13g2_decap_8 FILLER_35_855 ();
 sg13g2_decap_8 FILLER_35_862 ();
 sg13g2_decap_8 FILLER_35_869 ();
 sg13g2_decap_8 FILLER_35_876 ();
 sg13g2_decap_8 FILLER_35_883 ();
 sg13g2_decap_8 FILLER_35_890 ();
 sg13g2_decap_8 FILLER_35_897 ();
 sg13g2_decap_8 FILLER_35_904 ();
 sg13g2_decap_8 FILLER_35_911 ();
 sg13g2_decap_8 FILLER_35_918 ();
 sg13g2_decap_8 FILLER_35_925 ();
 sg13g2_decap_8 FILLER_35_932 ();
 sg13g2_decap_8 FILLER_35_939 ();
 sg13g2_decap_8 FILLER_35_946 ();
 sg13g2_decap_8 FILLER_35_953 ();
 sg13g2_decap_8 FILLER_35_960 ();
 sg13g2_decap_8 FILLER_35_967 ();
 sg13g2_decap_8 FILLER_35_974 ();
 sg13g2_decap_8 FILLER_35_981 ();
 sg13g2_decap_8 FILLER_35_988 ();
 sg13g2_decap_8 FILLER_35_995 ();
 sg13g2_decap_8 FILLER_35_1002 ();
 sg13g2_decap_8 FILLER_35_1009 ();
 sg13g2_decap_8 FILLER_35_1016 ();
 sg13g2_decap_4 FILLER_35_1023 ();
 sg13g2_fill_2 FILLER_35_1027 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_34 ();
 sg13g2_fill_1 FILLER_36_81 ();
 sg13g2_fill_2 FILLER_36_95 ();
 sg13g2_fill_1 FILLER_36_97 ();
 sg13g2_decap_8 FILLER_36_101 ();
 sg13g2_decap_4 FILLER_36_108 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_decap_4 FILLER_36_165 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_decap_4 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_decap_4 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_decap_4 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_decap_8 FILLER_36_298 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_4 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_fill_2 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_fill_1 FILLER_36_379 ();
 sg13g2_decap_4 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_decap_4 FILLER_36_471 ();
 sg13g2_fill_2 FILLER_36_475 ();
 sg13g2_decap_8 FILLER_36_531 ();
 sg13g2_decap_8 FILLER_36_538 ();
 sg13g2_decap_8 FILLER_36_545 ();
 sg13g2_decap_8 FILLER_36_552 ();
 sg13g2_decap_8 FILLER_36_559 ();
 sg13g2_decap_8 FILLER_36_566 ();
 sg13g2_decap_8 FILLER_36_573 ();
 sg13g2_decap_8 FILLER_36_580 ();
 sg13g2_decap_8 FILLER_36_587 ();
 sg13g2_decap_8 FILLER_36_594 ();
 sg13g2_decap_8 FILLER_36_601 ();
 sg13g2_decap_8 FILLER_36_608 ();
 sg13g2_decap_8 FILLER_36_615 ();
 sg13g2_decap_8 FILLER_36_622 ();
 sg13g2_decap_8 FILLER_36_629 ();
 sg13g2_decap_8 FILLER_36_636 ();
 sg13g2_decap_8 FILLER_36_643 ();
 sg13g2_decap_8 FILLER_36_650 ();
 sg13g2_decap_8 FILLER_36_657 ();
 sg13g2_decap_8 FILLER_36_664 ();
 sg13g2_decap_8 FILLER_36_671 ();
 sg13g2_decap_8 FILLER_36_678 ();
 sg13g2_decap_8 FILLER_36_685 ();
 sg13g2_decap_8 FILLER_36_692 ();
 sg13g2_decap_8 FILLER_36_699 ();
 sg13g2_decap_8 FILLER_36_706 ();
 sg13g2_decap_8 FILLER_36_713 ();
 sg13g2_decap_8 FILLER_36_720 ();
 sg13g2_decap_8 FILLER_36_727 ();
 sg13g2_decap_8 FILLER_36_734 ();
 sg13g2_decap_8 FILLER_36_741 ();
 sg13g2_decap_8 FILLER_36_748 ();
 sg13g2_decap_8 FILLER_36_755 ();
 sg13g2_decap_8 FILLER_36_762 ();
 sg13g2_decap_8 FILLER_36_769 ();
 sg13g2_decap_8 FILLER_36_776 ();
 sg13g2_decap_8 FILLER_36_783 ();
 sg13g2_decap_8 FILLER_36_790 ();
 sg13g2_decap_8 FILLER_36_797 ();
 sg13g2_decap_8 FILLER_36_804 ();
 sg13g2_decap_8 FILLER_36_811 ();
 sg13g2_decap_8 FILLER_36_818 ();
 sg13g2_decap_8 FILLER_36_825 ();
 sg13g2_decap_8 FILLER_36_832 ();
 sg13g2_decap_8 FILLER_36_839 ();
 sg13g2_decap_8 FILLER_36_846 ();
 sg13g2_decap_8 FILLER_36_853 ();
 sg13g2_decap_8 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_36_867 ();
 sg13g2_decap_8 FILLER_36_874 ();
 sg13g2_decap_8 FILLER_36_881 ();
 sg13g2_decap_8 FILLER_36_888 ();
 sg13g2_decap_8 FILLER_36_895 ();
 sg13g2_decap_8 FILLER_36_902 ();
 sg13g2_decap_8 FILLER_36_909 ();
 sg13g2_decap_8 FILLER_36_916 ();
 sg13g2_decap_8 FILLER_36_923 ();
 sg13g2_decap_8 FILLER_36_930 ();
 sg13g2_decap_8 FILLER_36_937 ();
 sg13g2_decap_8 FILLER_36_944 ();
 sg13g2_decap_8 FILLER_36_951 ();
 sg13g2_decap_8 FILLER_36_958 ();
 sg13g2_decap_8 FILLER_36_965 ();
 sg13g2_decap_8 FILLER_36_972 ();
 sg13g2_decap_8 FILLER_36_979 ();
 sg13g2_decap_8 FILLER_36_986 ();
 sg13g2_decap_8 FILLER_36_993 ();
 sg13g2_decap_8 FILLER_36_1000 ();
 sg13g2_decap_8 FILLER_36_1007 ();
 sg13g2_decap_8 FILLER_36_1014 ();
 sg13g2_decap_8 FILLER_36_1021 ();
 sg13g2_fill_1 FILLER_36_1028 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_11 ();
 sg13g2_decap_4 FILLER_37_16 ();
 sg13g2_fill_2 FILLER_37_20 ();
 sg13g2_fill_1 FILLER_37_45 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_fill_1 FILLER_37_106 ();
 sg13g2_decap_4 FILLER_37_134 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_163 ();
 sg13g2_decap_8 FILLER_37_234 ();
 sg13g2_decap_8 FILLER_37_241 ();
 sg13g2_decap_8 FILLER_37_248 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_282 ();
 sg13g2_decap_4 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_fill_2 FILLER_37_395 ();
 sg13g2_fill_1 FILLER_37_397 ();
 sg13g2_decap_8 FILLER_37_411 ();
 sg13g2_fill_1 FILLER_37_418 ();
 sg13g2_decap_8 FILLER_37_473 ();
 sg13g2_fill_2 FILLER_37_480 ();
 sg13g2_fill_1 FILLER_37_482 ();
 sg13g2_fill_1 FILLER_37_496 ();
 sg13g2_decap_8 FILLER_37_533 ();
 sg13g2_decap_8 FILLER_37_540 ();
 sg13g2_decap_8 FILLER_37_547 ();
 sg13g2_decap_8 FILLER_37_554 ();
 sg13g2_decap_8 FILLER_37_561 ();
 sg13g2_decap_8 FILLER_37_568 ();
 sg13g2_decap_8 FILLER_37_575 ();
 sg13g2_decap_8 FILLER_37_582 ();
 sg13g2_decap_8 FILLER_37_589 ();
 sg13g2_decap_8 FILLER_37_596 ();
 sg13g2_decap_8 FILLER_37_603 ();
 sg13g2_decap_8 FILLER_37_610 ();
 sg13g2_decap_8 FILLER_37_617 ();
 sg13g2_decap_8 FILLER_37_624 ();
 sg13g2_decap_8 FILLER_37_631 ();
 sg13g2_decap_8 FILLER_37_638 ();
 sg13g2_decap_8 FILLER_37_645 ();
 sg13g2_decap_8 FILLER_37_652 ();
 sg13g2_decap_8 FILLER_37_659 ();
 sg13g2_decap_8 FILLER_37_666 ();
 sg13g2_decap_8 FILLER_37_673 ();
 sg13g2_decap_8 FILLER_37_680 ();
 sg13g2_decap_8 FILLER_37_687 ();
 sg13g2_decap_8 FILLER_37_694 ();
 sg13g2_decap_8 FILLER_37_701 ();
 sg13g2_decap_8 FILLER_37_708 ();
 sg13g2_decap_8 FILLER_37_715 ();
 sg13g2_decap_8 FILLER_37_722 ();
 sg13g2_decap_8 FILLER_37_729 ();
 sg13g2_decap_8 FILLER_37_736 ();
 sg13g2_decap_8 FILLER_37_743 ();
 sg13g2_decap_8 FILLER_37_750 ();
 sg13g2_decap_8 FILLER_37_757 ();
 sg13g2_decap_8 FILLER_37_764 ();
 sg13g2_decap_8 FILLER_37_771 ();
 sg13g2_decap_8 FILLER_37_778 ();
 sg13g2_decap_8 FILLER_37_785 ();
 sg13g2_decap_8 FILLER_37_792 ();
 sg13g2_decap_8 FILLER_37_799 ();
 sg13g2_decap_8 FILLER_37_806 ();
 sg13g2_decap_8 FILLER_37_813 ();
 sg13g2_decap_8 FILLER_37_820 ();
 sg13g2_decap_8 FILLER_37_827 ();
 sg13g2_decap_8 FILLER_37_834 ();
 sg13g2_decap_8 FILLER_37_841 ();
 sg13g2_decap_8 FILLER_37_848 ();
 sg13g2_decap_8 FILLER_37_855 ();
 sg13g2_decap_8 FILLER_37_862 ();
 sg13g2_decap_8 FILLER_37_869 ();
 sg13g2_decap_8 FILLER_37_876 ();
 sg13g2_decap_8 FILLER_37_883 ();
 sg13g2_decap_8 FILLER_37_890 ();
 sg13g2_decap_8 FILLER_37_897 ();
 sg13g2_decap_8 FILLER_37_904 ();
 sg13g2_decap_8 FILLER_37_911 ();
 sg13g2_decap_8 FILLER_37_918 ();
 sg13g2_decap_8 FILLER_37_925 ();
 sg13g2_decap_8 FILLER_37_932 ();
 sg13g2_decap_8 FILLER_37_939 ();
 sg13g2_decap_8 FILLER_37_946 ();
 sg13g2_decap_8 FILLER_37_953 ();
 sg13g2_decap_8 FILLER_37_960 ();
 sg13g2_decap_8 FILLER_37_967 ();
 sg13g2_decap_8 FILLER_37_974 ();
 sg13g2_decap_8 FILLER_37_981 ();
 sg13g2_decap_8 FILLER_37_988 ();
 sg13g2_decap_8 FILLER_37_995 ();
 sg13g2_decap_8 FILLER_37_1002 ();
 sg13g2_decap_8 FILLER_37_1009 ();
 sg13g2_decap_8 FILLER_37_1016 ();
 sg13g2_decap_4 FILLER_37_1023 ();
 sg13g2_fill_2 FILLER_37_1027 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_33 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_113 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_decap_8 FILLER_38_176 ();
 sg13g2_decap_4 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_382 ();
 sg13g2_decap_4 FILLER_38_388 ();
 sg13g2_fill_2 FILLER_38_493 ();
 sg13g2_decap_8 FILLER_38_522 ();
 sg13g2_decap_8 FILLER_38_529 ();
 sg13g2_decap_8 FILLER_38_536 ();
 sg13g2_decap_8 FILLER_38_543 ();
 sg13g2_decap_8 FILLER_38_550 ();
 sg13g2_decap_8 FILLER_38_557 ();
 sg13g2_decap_8 FILLER_38_564 ();
 sg13g2_decap_8 FILLER_38_571 ();
 sg13g2_decap_8 FILLER_38_578 ();
 sg13g2_decap_8 FILLER_38_585 ();
 sg13g2_decap_8 FILLER_38_592 ();
 sg13g2_decap_8 FILLER_38_599 ();
 sg13g2_decap_8 FILLER_38_606 ();
 sg13g2_decap_8 FILLER_38_613 ();
 sg13g2_decap_8 FILLER_38_620 ();
 sg13g2_decap_8 FILLER_38_627 ();
 sg13g2_decap_8 FILLER_38_634 ();
 sg13g2_decap_8 FILLER_38_641 ();
 sg13g2_decap_8 FILLER_38_648 ();
 sg13g2_decap_8 FILLER_38_655 ();
 sg13g2_decap_8 FILLER_38_662 ();
 sg13g2_decap_8 FILLER_38_669 ();
 sg13g2_decap_8 FILLER_38_676 ();
 sg13g2_decap_8 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_690 ();
 sg13g2_decap_8 FILLER_38_697 ();
 sg13g2_decap_8 FILLER_38_704 ();
 sg13g2_decap_8 FILLER_38_711 ();
 sg13g2_decap_8 FILLER_38_718 ();
 sg13g2_decap_8 FILLER_38_725 ();
 sg13g2_decap_8 FILLER_38_732 ();
 sg13g2_decap_8 FILLER_38_739 ();
 sg13g2_decap_8 FILLER_38_746 ();
 sg13g2_decap_8 FILLER_38_753 ();
 sg13g2_decap_8 FILLER_38_760 ();
 sg13g2_decap_8 FILLER_38_767 ();
 sg13g2_decap_8 FILLER_38_774 ();
 sg13g2_decap_8 FILLER_38_781 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_decap_8 FILLER_38_795 ();
 sg13g2_decap_8 FILLER_38_802 ();
 sg13g2_decap_8 FILLER_38_809 ();
 sg13g2_decap_8 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_830 ();
 sg13g2_decap_8 FILLER_38_837 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_8 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_38_865 ();
 sg13g2_decap_8 FILLER_38_872 ();
 sg13g2_decap_8 FILLER_38_879 ();
 sg13g2_decap_8 FILLER_38_886 ();
 sg13g2_decap_8 FILLER_38_893 ();
 sg13g2_decap_8 FILLER_38_900 ();
 sg13g2_decap_8 FILLER_38_907 ();
 sg13g2_decap_8 FILLER_38_914 ();
 sg13g2_decap_8 FILLER_38_921 ();
 sg13g2_decap_8 FILLER_38_928 ();
 sg13g2_decap_8 FILLER_38_935 ();
 sg13g2_decap_8 FILLER_38_942 ();
 sg13g2_decap_8 FILLER_38_949 ();
 sg13g2_decap_8 FILLER_38_956 ();
 sg13g2_decap_8 FILLER_38_963 ();
 sg13g2_decap_8 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_8 FILLER_38_991 ();
 sg13g2_decap_8 FILLER_38_998 ();
 sg13g2_decap_8 FILLER_38_1005 ();
 sg13g2_decap_8 FILLER_38_1012 ();
 sg13g2_decap_8 FILLER_38_1019 ();
 sg13g2_fill_2 FILLER_38_1026 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_34 ();
 sg13g2_fill_2 FILLER_39_53 ();
 sg13g2_fill_2 FILLER_39_85 ();
 sg13g2_decap_8 FILLER_39_100 ();
 sg13g2_decap_8 FILLER_39_165 ();
 sg13g2_fill_2 FILLER_39_172 ();
 sg13g2_fill_1 FILLER_39_174 ();
 sg13g2_decap_8 FILLER_39_179 ();
 sg13g2_fill_2 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_256 ();
 sg13g2_fill_1 FILLER_39_258 ();
 sg13g2_fill_2 FILLER_39_287 ();
 sg13g2_fill_2 FILLER_39_294 ();
 sg13g2_fill_1 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_366 ();
 sg13g2_fill_2 FILLER_39_377 ();
 sg13g2_decap_8 FILLER_39_383 ();
 sg13g2_fill_1 FILLER_39_432 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_fill_1 FILLER_39_476 ();
 sg13g2_fill_2 FILLER_39_488 ();
 sg13g2_fill_1 FILLER_39_495 ();
 sg13g2_fill_2 FILLER_39_501 ();
 sg13g2_decap_8 FILLER_39_520 ();
 sg13g2_decap_8 FILLER_39_527 ();
 sg13g2_decap_8 FILLER_39_534 ();
 sg13g2_decap_8 FILLER_39_541 ();
 sg13g2_decap_8 FILLER_39_548 ();
 sg13g2_decap_8 FILLER_39_555 ();
 sg13g2_decap_8 FILLER_39_562 ();
 sg13g2_decap_8 FILLER_39_569 ();
 sg13g2_decap_8 FILLER_39_576 ();
 sg13g2_decap_8 FILLER_39_583 ();
 sg13g2_decap_8 FILLER_39_590 ();
 sg13g2_decap_8 FILLER_39_597 ();
 sg13g2_decap_8 FILLER_39_604 ();
 sg13g2_decap_8 FILLER_39_611 ();
 sg13g2_decap_8 FILLER_39_618 ();
 sg13g2_decap_8 FILLER_39_625 ();
 sg13g2_decap_8 FILLER_39_632 ();
 sg13g2_decap_8 FILLER_39_639 ();
 sg13g2_decap_8 FILLER_39_646 ();
 sg13g2_decap_8 FILLER_39_653 ();
 sg13g2_decap_8 FILLER_39_660 ();
 sg13g2_decap_8 FILLER_39_667 ();
 sg13g2_decap_8 FILLER_39_674 ();
 sg13g2_decap_8 FILLER_39_681 ();
 sg13g2_decap_8 FILLER_39_688 ();
 sg13g2_decap_8 FILLER_39_695 ();
 sg13g2_decap_8 FILLER_39_702 ();
 sg13g2_decap_8 FILLER_39_709 ();
 sg13g2_decap_8 FILLER_39_716 ();
 sg13g2_decap_8 FILLER_39_723 ();
 sg13g2_decap_8 FILLER_39_730 ();
 sg13g2_decap_8 FILLER_39_737 ();
 sg13g2_decap_8 FILLER_39_744 ();
 sg13g2_decap_8 FILLER_39_751 ();
 sg13g2_decap_8 FILLER_39_758 ();
 sg13g2_decap_8 FILLER_39_765 ();
 sg13g2_decap_8 FILLER_39_772 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_decap_8 FILLER_39_814 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_8 FILLER_39_856 ();
 sg13g2_decap_8 FILLER_39_863 ();
 sg13g2_decap_8 FILLER_39_870 ();
 sg13g2_decap_8 FILLER_39_877 ();
 sg13g2_decap_8 FILLER_39_884 ();
 sg13g2_decap_8 FILLER_39_891 ();
 sg13g2_decap_8 FILLER_39_898 ();
 sg13g2_decap_8 FILLER_39_905 ();
 sg13g2_decap_8 FILLER_39_912 ();
 sg13g2_decap_8 FILLER_39_919 ();
 sg13g2_decap_8 FILLER_39_926 ();
 sg13g2_decap_8 FILLER_39_933 ();
 sg13g2_decap_8 FILLER_39_940 ();
 sg13g2_decap_8 FILLER_39_947 ();
 sg13g2_decap_8 FILLER_39_954 ();
 sg13g2_decap_8 FILLER_39_961 ();
 sg13g2_decap_8 FILLER_39_968 ();
 sg13g2_decap_8 FILLER_39_975 ();
 sg13g2_decap_8 FILLER_39_982 ();
 sg13g2_decap_8 FILLER_39_989 ();
 sg13g2_decap_8 FILLER_39_996 ();
 sg13g2_decap_8 FILLER_39_1003 ();
 sg13g2_decap_8 FILLER_39_1010 ();
 sg13g2_decap_8 FILLER_39_1017 ();
 sg13g2_decap_4 FILLER_39_1024 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_7 ();
 sg13g2_fill_2 FILLER_40_11 ();
 sg13g2_decap_8 FILLER_40_17 ();
 sg13g2_decap_4 FILLER_40_24 ();
 sg13g2_fill_1 FILLER_40_28 ();
 sg13g2_fill_2 FILLER_40_53 ();
 sg13g2_fill_1 FILLER_40_96 ();
 sg13g2_fill_2 FILLER_40_150 ();
 sg13g2_fill_1 FILLER_40_164 ();
 sg13g2_decap_8 FILLER_40_218 ();
 sg13g2_decap_4 FILLER_40_225 ();
 sg13g2_fill_2 FILLER_40_229 ();
 sg13g2_decap_8 FILLER_40_235 ();
 sg13g2_fill_2 FILLER_40_242 ();
 sg13g2_fill_2 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_262 ();
 sg13g2_fill_1 FILLER_40_277 ();
 sg13g2_fill_2 FILLER_40_334 ();
 sg13g2_fill_2 FILLER_40_355 ();
 sg13g2_fill_1 FILLER_40_357 ();
 sg13g2_decap_4 FILLER_40_385 ();
 sg13g2_fill_1 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_513 ();
 sg13g2_decap_8 FILLER_40_520 ();
 sg13g2_decap_8 FILLER_40_527 ();
 sg13g2_decap_8 FILLER_40_534 ();
 sg13g2_decap_8 FILLER_40_541 ();
 sg13g2_decap_8 FILLER_40_548 ();
 sg13g2_decap_8 FILLER_40_555 ();
 sg13g2_decap_8 FILLER_40_562 ();
 sg13g2_decap_8 FILLER_40_569 ();
 sg13g2_decap_8 FILLER_40_576 ();
 sg13g2_decap_8 FILLER_40_583 ();
 sg13g2_decap_8 FILLER_40_590 ();
 sg13g2_decap_8 FILLER_40_597 ();
 sg13g2_decap_8 FILLER_40_604 ();
 sg13g2_decap_8 FILLER_40_611 ();
 sg13g2_decap_8 FILLER_40_618 ();
 sg13g2_decap_8 FILLER_40_625 ();
 sg13g2_decap_8 FILLER_40_632 ();
 sg13g2_decap_8 FILLER_40_639 ();
 sg13g2_decap_8 FILLER_40_646 ();
 sg13g2_decap_8 FILLER_40_653 ();
 sg13g2_decap_8 FILLER_40_660 ();
 sg13g2_decap_8 FILLER_40_667 ();
 sg13g2_decap_8 FILLER_40_674 ();
 sg13g2_decap_8 FILLER_40_681 ();
 sg13g2_decap_8 FILLER_40_688 ();
 sg13g2_decap_8 FILLER_40_695 ();
 sg13g2_decap_8 FILLER_40_702 ();
 sg13g2_decap_8 FILLER_40_709 ();
 sg13g2_decap_8 FILLER_40_716 ();
 sg13g2_decap_8 FILLER_40_723 ();
 sg13g2_decap_8 FILLER_40_730 ();
 sg13g2_decap_8 FILLER_40_737 ();
 sg13g2_decap_8 FILLER_40_744 ();
 sg13g2_decap_8 FILLER_40_751 ();
 sg13g2_decap_8 FILLER_40_758 ();
 sg13g2_decap_8 FILLER_40_765 ();
 sg13g2_decap_8 FILLER_40_772 ();
 sg13g2_decap_8 FILLER_40_779 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_800 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_828 ();
 sg13g2_decap_8 FILLER_40_835 ();
 sg13g2_decap_8 FILLER_40_842 ();
 sg13g2_decap_8 FILLER_40_849 ();
 sg13g2_decap_8 FILLER_40_856 ();
 sg13g2_decap_8 FILLER_40_863 ();
 sg13g2_decap_8 FILLER_40_870 ();
 sg13g2_decap_8 FILLER_40_877 ();
 sg13g2_decap_8 FILLER_40_884 ();
 sg13g2_decap_8 FILLER_40_891 ();
 sg13g2_decap_8 FILLER_40_898 ();
 sg13g2_decap_8 FILLER_40_905 ();
 sg13g2_decap_8 FILLER_40_912 ();
 sg13g2_decap_8 FILLER_40_919 ();
 sg13g2_decap_8 FILLER_40_926 ();
 sg13g2_decap_8 FILLER_40_933 ();
 sg13g2_decap_8 FILLER_40_940 ();
 sg13g2_decap_8 FILLER_40_947 ();
 sg13g2_decap_8 FILLER_40_954 ();
 sg13g2_decap_8 FILLER_40_961 ();
 sg13g2_decap_8 FILLER_40_968 ();
 sg13g2_decap_8 FILLER_40_975 ();
 sg13g2_decap_8 FILLER_40_982 ();
 sg13g2_decap_8 FILLER_40_989 ();
 sg13g2_decap_8 FILLER_40_996 ();
 sg13g2_decap_8 FILLER_40_1003 ();
 sg13g2_decap_8 FILLER_40_1010 ();
 sg13g2_decap_8 FILLER_40_1017 ();
 sg13g2_decap_4 FILLER_40_1024 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_34 ();
 sg13g2_fill_1 FILLER_41_75 ();
 sg13g2_fill_1 FILLER_41_179 ();
 sg13g2_decap_8 FILLER_41_230 ();
 sg13g2_fill_1 FILLER_41_237 ();
 sg13g2_decap_8 FILLER_41_243 ();
 sg13g2_fill_2 FILLER_41_250 ();
 sg13g2_fill_1 FILLER_41_324 ();
 sg13g2_fill_2 FILLER_41_371 ();
 sg13g2_fill_1 FILLER_41_373 ();
 sg13g2_decap_8 FILLER_41_377 ();
 sg13g2_fill_1 FILLER_41_384 ();
 sg13g2_fill_1 FILLER_41_397 ();
 sg13g2_fill_2 FILLER_41_427 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_fill_1 FILLER_41_458 ();
 sg13g2_fill_1 FILLER_41_486 ();
 sg13g2_decap_4 FILLER_41_501 ();
 sg13g2_decap_8 FILLER_41_514 ();
 sg13g2_decap_8 FILLER_41_521 ();
 sg13g2_decap_8 FILLER_41_528 ();
 sg13g2_decap_8 FILLER_41_535 ();
 sg13g2_decap_8 FILLER_41_542 ();
 sg13g2_decap_8 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_556 ();
 sg13g2_decap_8 FILLER_41_563 ();
 sg13g2_decap_8 FILLER_41_570 ();
 sg13g2_decap_8 FILLER_41_577 ();
 sg13g2_decap_8 FILLER_41_584 ();
 sg13g2_decap_8 FILLER_41_591 ();
 sg13g2_decap_8 FILLER_41_598 ();
 sg13g2_decap_8 FILLER_41_605 ();
 sg13g2_decap_8 FILLER_41_612 ();
 sg13g2_decap_8 FILLER_41_619 ();
 sg13g2_decap_8 FILLER_41_626 ();
 sg13g2_decap_8 FILLER_41_633 ();
 sg13g2_decap_8 FILLER_41_640 ();
 sg13g2_decap_8 FILLER_41_647 ();
 sg13g2_decap_8 FILLER_41_654 ();
 sg13g2_decap_8 FILLER_41_661 ();
 sg13g2_decap_8 FILLER_41_668 ();
 sg13g2_decap_8 FILLER_41_675 ();
 sg13g2_decap_8 FILLER_41_682 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_710 ();
 sg13g2_decap_8 FILLER_41_717 ();
 sg13g2_decap_8 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_731 ();
 sg13g2_decap_8 FILLER_41_738 ();
 sg13g2_decap_8 FILLER_41_745 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_773 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_794 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_8 FILLER_41_857 ();
 sg13g2_decap_8 FILLER_41_864 ();
 sg13g2_decap_8 FILLER_41_871 ();
 sg13g2_decap_8 FILLER_41_878 ();
 sg13g2_decap_8 FILLER_41_885 ();
 sg13g2_decap_8 FILLER_41_892 ();
 sg13g2_decap_8 FILLER_41_899 ();
 sg13g2_decap_8 FILLER_41_906 ();
 sg13g2_decap_8 FILLER_41_913 ();
 sg13g2_decap_8 FILLER_41_920 ();
 sg13g2_decap_8 FILLER_41_927 ();
 sg13g2_decap_8 FILLER_41_934 ();
 sg13g2_decap_8 FILLER_41_941 ();
 sg13g2_decap_8 FILLER_41_948 ();
 sg13g2_decap_8 FILLER_41_955 ();
 sg13g2_decap_8 FILLER_41_962 ();
 sg13g2_decap_8 FILLER_41_969 ();
 sg13g2_decap_8 FILLER_41_976 ();
 sg13g2_decap_8 FILLER_41_983 ();
 sg13g2_decap_8 FILLER_41_990 ();
 sg13g2_decap_8 FILLER_41_997 ();
 sg13g2_decap_8 FILLER_41_1004 ();
 sg13g2_decap_8 FILLER_41_1011 ();
 sg13g2_decap_8 FILLER_41_1018 ();
 sg13g2_decap_4 FILLER_41_1025 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_4 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_34 ();
 sg13g2_fill_1 FILLER_42_58 ();
 sg13g2_fill_2 FILLER_42_105 ();
 sg13g2_fill_1 FILLER_42_107 ();
 sg13g2_decap_8 FILLER_42_218 ();
 sg13g2_decap_8 FILLER_42_225 ();
 sg13g2_decap_4 FILLER_42_232 ();
 sg13g2_fill_2 FILLER_42_294 ();
 sg13g2_fill_1 FILLER_42_344 ();
 sg13g2_decap_8 FILLER_42_358 ();
 sg13g2_decap_4 FILLER_42_365 ();
 sg13g2_fill_2 FILLER_42_455 ();
 sg13g2_fill_1 FILLER_42_457 ();
 sg13g2_decap_8 FILLER_42_471 ();
 sg13g2_decap_4 FILLER_42_478 ();
 sg13g2_fill_1 FILLER_42_482 ();
 sg13g2_decap_8 FILLER_42_496 ();
 sg13g2_decap_8 FILLER_42_503 ();
 sg13g2_decap_8 FILLER_42_510 ();
 sg13g2_decap_8 FILLER_42_517 ();
 sg13g2_decap_8 FILLER_42_524 ();
 sg13g2_decap_8 FILLER_42_531 ();
 sg13g2_decap_8 FILLER_42_538 ();
 sg13g2_decap_8 FILLER_42_545 ();
 sg13g2_decap_8 FILLER_42_552 ();
 sg13g2_decap_8 FILLER_42_559 ();
 sg13g2_decap_8 FILLER_42_566 ();
 sg13g2_decap_8 FILLER_42_573 ();
 sg13g2_decap_8 FILLER_42_580 ();
 sg13g2_decap_8 FILLER_42_587 ();
 sg13g2_decap_8 FILLER_42_594 ();
 sg13g2_decap_8 FILLER_42_601 ();
 sg13g2_decap_8 FILLER_42_608 ();
 sg13g2_decap_8 FILLER_42_615 ();
 sg13g2_decap_8 FILLER_42_622 ();
 sg13g2_decap_8 FILLER_42_629 ();
 sg13g2_decap_8 FILLER_42_636 ();
 sg13g2_decap_8 FILLER_42_643 ();
 sg13g2_decap_8 FILLER_42_650 ();
 sg13g2_decap_8 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_664 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_decap_8 FILLER_42_678 ();
 sg13g2_decap_8 FILLER_42_685 ();
 sg13g2_decap_8 FILLER_42_692 ();
 sg13g2_decap_8 FILLER_42_699 ();
 sg13g2_decap_8 FILLER_42_706 ();
 sg13g2_decap_8 FILLER_42_713 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_decap_8 FILLER_42_727 ();
 sg13g2_decap_8 FILLER_42_734 ();
 sg13g2_decap_8 FILLER_42_741 ();
 sg13g2_decap_8 FILLER_42_748 ();
 sg13g2_decap_8 FILLER_42_755 ();
 sg13g2_decap_8 FILLER_42_762 ();
 sg13g2_decap_8 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_776 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_decap_8 FILLER_42_790 ();
 sg13g2_decap_8 FILLER_42_797 ();
 sg13g2_decap_8 FILLER_42_804 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_decap_8 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_42_867 ();
 sg13g2_decap_8 FILLER_42_874 ();
 sg13g2_decap_8 FILLER_42_881 ();
 sg13g2_decap_8 FILLER_42_888 ();
 sg13g2_decap_8 FILLER_42_895 ();
 sg13g2_decap_8 FILLER_42_902 ();
 sg13g2_decap_8 FILLER_42_909 ();
 sg13g2_decap_8 FILLER_42_916 ();
 sg13g2_decap_8 FILLER_42_923 ();
 sg13g2_decap_8 FILLER_42_930 ();
 sg13g2_decap_8 FILLER_42_937 ();
 sg13g2_decap_8 FILLER_42_944 ();
 sg13g2_decap_8 FILLER_42_951 ();
 sg13g2_decap_8 FILLER_42_958 ();
 sg13g2_decap_8 FILLER_42_965 ();
 sg13g2_decap_8 FILLER_42_972 ();
 sg13g2_decap_8 FILLER_42_979 ();
 sg13g2_decap_8 FILLER_42_986 ();
 sg13g2_decap_8 FILLER_42_993 ();
 sg13g2_decap_8 FILLER_42_1000 ();
 sg13g2_decap_8 FILLER_42_1007 ();
 sg13g2_decap_8 FILLER_42_1014 ();
 sg13g2_decap_8 FILLER_42_1021 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_58 ();
 sg13g2_fill_1 FILLER_43_64 ();
 sg13g2_decap_4 FILLER_43_78 ();
 sg13g2_decap_4 FILLER_43_96 ();
 sg13g2_fill_2 FILLER_43_100 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_4 FILLER_43_168 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_2 FILLER_43_184 ();
 sg13g2_fill_1 FILLER_43_186 ();
 sg13g2_fill_2 FILLER_43_208 ();
 sg13g2_decap_8 FILLER_43_223 ();
 sg13g2_decap_8 FILLER_43_230 ();
 sg13g2_fill_1 FILLER_43_237 ();
 sg13g2_fill_2 FILLER_43_251 ();
 sg13g2_fill_1 FILLER_43_253 ();
 sg13g2_fill_1 FILLER_43_258 ();
 sg13g2_fill_2 FILLER_43_269 ();
 sg13g2_fill_1 FILLER_43_271 ();
 sg13g2_fill_1 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_365 ();
 sg13g2_fill_2 FILLER_43_386 ();
 sg13g2_fill_1 FILLER_43_388 ();
 sg13g2_fill_2 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_474 ();
 sg13g2_decap_8 FILLER_43_481 ();
 sg13g2_decap_8 FILLER_43_488 ();
 sg13g2_decap_8 FILLER_43_495 ();
 sg13g2_decap_8 FILLER_43_502 ();
 sg13g2_decap_8 FILLER_43_509 ();
 sg13g2_decap_8 FILLER_43_516 ();
 sg13g2_decap_8 FILLER_43_523 ();
 sg13g2_decap_8 FILLER_43_530 ();
 sg13g2_decap_8 FILLER_43_537 ();
 sg13g2_decap_8 FILLER_43_544 ();
 sg13g2_decap_8 FILLER_43_551 ();
 sg13g2_decap_8 FILLER_43_558 ();
 sg13g2_decap_8 FILLER_43_565 ();
 sg13g2_decap_8 FILLER_43_572 ();
 sg13g2_decap_8 FILLER_43_579 ();
 sg13g2_decap_8 FILLER_43_586 ();
 sg13g2_decap_8 FILLER_43_593 ();
 sg13g2_decap_8 FILLER_43_600 ();
 sg13g2_decap_8 FILLER_43_607 ();
 sg13g2_decap_8 FILLER_43_614 ();
 sg13g2_decap_8 FILLER_43_621 ();
 sg13g2_decap_8 FILLER_43_628 ();
 sg13g2_decap_8 FILLER_43_635 ();
 sg13g2_decap_8 FILLER_43_642 ();
 sg13g2_decap_8 FILLER_43_649 ();
 sg13g2_decap_8 FILLER_43_656 ();
 sg13g2_decap_8 FILLER_43_663 ();
 sg13g2_decap_8 FILLER_43_670 ();
 sg13g2_decap_8 FILLER_43_677 ();
 sg13g2_decap_8 FILLER_43_684 ();
 sg13g2_decap_8 FILLER_43_691 ();
 sg13g2_decap_8 FILLER_43_698 ();
 sg13g2_decap_8 FILLER_43_705 ();
 sg13g2_decap_8 FILLER_43_712 ();
 sg13g2_decap_8 FILLER_43_719 ();
 sg13g2_decap_8 FILLER_43_726 ();
 sg13g2_decap_8 FILLER_43_733 ();
 sg13g2_decap_8 FILLER_43_740 ();
 sg13g2_decap_8 FILLER_43_747 ();
 sg13g2_decap_8 FILLER_43_754 ();
 sg13g2_decap_8 FILLER_43_761 ();
 sg13g2_decap_8 FILLER_43_768 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_782 ();
 sg13g2_decap_8 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_796 ();
 sg13g2_decap_8 FILLER_43_803 ();
 sg13g2_decap_8 FILLER_43_810 ();
 sg13g2_decap_8 FILLER_43_817 ();
 sg13g2_decap_8 FILLER_43_824 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_8 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_decap_8 FILLER_43_859 ();
 sg13g2_decap_8 FILLER_43_866 ();
 sg13g2_decap_8 FILLER_43_873 ();
 sg13g2_decap_8 FILLER_43_880 ();
 sg13g2_decap_8 FILLER_43_887 ();
 sg13g2_decap_8 FILLER_43_894 ();
 sg13g2_decap_8 FILLER_43_901 ();
 sg13g2_decap_8 FILLER_43_908 ();
 sg13g2_decap_8 FILLER_43_915 ();
 sg13g2_decap_8 FILLER_43_922 ();
 sg13g2_decap_8 FILLER_43_929 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_decap_8 FILLER_43_950 ();
 sg13g2_decap_8 FILLER_43_957 ();
 sg13g2_decap_8 FILLER_43_964 ();
 sg13g2_decap_8 FILLER_43_971 ();
 sg13g2_decap_8 FILLER_43_978 ();
 sg13g2_decap_8 FILLER_43_985 ();
 sg13g2_decap_8 FILLER_43_992 ();
 sg13g2_decap_8 FILLER_43_999 ();
 sg13g2_decap_8 FILLER_43_1006 ();
 sg13g2_decap_8 FILLER_43_1013 ();
 sg13g2_decap_8 FILLER_43_1020 ();
 sg13g2_fill_2 FILLER_43_1027 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_4 FILLER_44_14 ();
 sg13g2_fill_2 FILLER_44_18 ();
 sg13g2_decap_8 FILLER_44_24 ();
 sg13g2_fill_1 FILLER_44_127 ();
 sg13g2_fill_1 FILLER_44_156 ();
 sg13g2_decap_8 FILLER_44_198 ();
 sg13g2_decap_8 FILLER_44_205 ();
 sg13g2_decap_4 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_243 ();
 sg13g2_fill_2 FILLER_44_256 ();
 sg13g2_fill_2 FILLER_44_276 ();
 sg13g2_fill_2 FILLER_44_302 ();
 sg13g2_fill_1 FILLER_44_322 ();
 sg13g2_fill_2 FILLER_44_395 ();
 sg13g2_fill_1 FILLER_44_397 ();
 sg13g2_fill_2 FILLER_44_444 ();
 sg13g2_decap_8 FILLER_44_459 ();
 sg13g2_decap_8 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_473 ();
 sg13g2_decap_8 FILLER_44_480 ();
 sg13g2_decap_8 FILLER_44_487 ();
 sg13g2_decap_8 FILLER_44_494 ();
 sg13g2_decap_8 FILLER_44_501 ();
 sg13g2_decap_8 FILLER_44_508 ();
 sg13g2_decap_8 FILLER_44_515 ();
 sg13g2_decap_8 FILLER_44_522 ();
 sg13g2_decap_8 FILLER_44_529 ();
 sg13g2_decap_8 FILLER_44_536 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_557 ();
 sg13g2_decap_8 FILLER_44_564 ();
 sg13g2_decap_8 FILLER_44_571 ();
 sg13g2_decap_8 FILLER_44_578 ();
 sg13g2_decap_8 FILLER_44_585 ();
 sg13g2_decap_8 FILLER_44_592 ();
 sg13g2_decap_8 FILLER_44_599 ();
 sg13g2_decap_8 FILLER_44_606 ();
 sg13g2_decap_8 FILLER_44_613 ();
 sg13g2_decap_8 FILLER_44_620 ();
 sg13g2_decap_8 FILLER_44_627 ();
 sg13g2_decap_8 FILLER_44_634 ();
 sg13g2_decap_8 FILLER_44_641 ();
 sg13g2_decap_8 FILLER_44_648 ();
 sg13g2_decap_8 FILLER_44_655 ();
 sg13g2_decap_8 FILLER_44_662 ();
 sg13g2_decap_8 FILLER_44_669 ();
 sg13g2_decap_8 FILLER_44_676 ();
 sg13g2_decap_8 FILLER_44_683 ();
 sg13g2_decap_8 FILLER_44_690 ();
 sg13g2_decap_8 FILLER_44_697 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_decap_8 FILLER_44_711 ();
 sg13g2_decap_8 FILLER_44_718 ();
 sg13g2_decap_8 FILLER_44_725 ();
 sg13g2_decap_8 FILLER_44_732 ();
 sg13g2_decap_8 FILLER_44_739 ();
 sg13g2_decap_8 FILLER_44_746 ();
 sg13g2_decap_8 FILLER_44_753 ();
 sg13g2_decap_8 FILLER_44_760 ();
 sg13g2_decap_8 FILLER_44_767 ();
 sg13g2_decap_8 FILLER_44_774 ();
 sg13g2_decap_8 FILLER_44_781 ();
 sg13g2_decap_8 FILLER_44_788 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_decap_8 FILLER_44_802 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_8 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_44_865 ();
 sg13g2_decap_8 FILLER_44_872 ();
 sg13g2_decap_8 FILLER_44_879 ();
 sg13g2_decap_8 FILLER_44_886 ();
 sg13g2_decap_8 FILLER_44_893 ();
 sg13g2_decap_8 FILLER_44_900 ();
 sg13g2_decap_8 FILLER_44_907 ();
 sg13g2_decap_8 FILLER_44_914 ();
 sg13g2_decap_8 FILLER_44_921 ();
 sg13g2_decap_8 FILLER_44_928 ();
 sg13g2_decap_8 FILLER_44_935 ();
 sg13g2_decap_8 FILLER_44_942 ();
 sg13g2_decap_8 FILLER_44_949 ();
 sg13g2_decap_8 FILLER_44_956 ();
 sg13g2_decap_8 FILLER_44_963 ();
 sg13g2_decap_8 FILLER_44_970 ();
 sg13g2_decap_8 FILLER_44_977 ();
 sg13g2_decap_8 FILLER_44_984 ();
 sg13g2_decap_8 FILLER_44_991 ();
 sg13g2_decap_8 FILLER_44_998 ();
 sg13g2_decap_8 FILLER_44_1005 ();
 sg13g2_decap_8 FILLER_44_1012 ();
 sg13g2_decap_8 FILLER_44_1019 ();
 sg13g2_fill_2 FILLER_44_1026 ();
 sg13g2_fill_1 FILLER_44_1028 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_35 ();
 sg13g2_fill_1 FILLER_45_39 ();
 sg13g2_decap_4 FILLER_45_44 ();
 sg13g2_fill_1 FILLER_45_48 ();
 sg13g2_fill_1 FILLER_45_72 ();
 sg13g2_fill_2 FILLER_45_82 ();
 sg13g2_fill_1 FILLER_45_84 ();
 sg13g2_decap_4 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_183 ();
 sg13g2_fill_2 FILLER_45_187 ();
 sg13g2_fill_2 FILLER_45_216 ();
 sg13g2_decap_4 FILLER_45_231 ();
 sg13g2_fill_2 FILLER_45_235 ();
 sg13g2_fill_2 FILLER_45_286 ();
 sg13g2_fill_1 FILLER_45_300 ();
 sg13g2_fill_2 FILLER_45_398 ();
 sg13g2_fill_2 FILLER_45_408 ();
 sg13g2_fill_1 FILLER_45_410 ();
 sg13g2_fill_2 FILLER_45_447 ();
 sg13g2_decap_8 FILLER_45_458 ();
 sg13g2_decap_8 FILLER_45_465 ();
 sg13g2_decap_8 FILLER_45_472 ();
 sg13g2_decap_8 FILLER_45_479 ();
 sg13g2_decap_8 FILLER_45_486 ();
 sg13g2_decap_8 FILLER_45_493 ();
 sg13g2_decap_8 FILLER_45_500 ();
 sg13g2_decap_8 FILLER_45_507 ();
 sg13g2_decap_8 FILLER_45_514 ();
 sg13g2_decap_8 FILLER_45_521 ();
 sg13g2_decap_8 FILLER_45_528 ();
 sg13g2_decap_8 FILLER_45_535 ();
 sg13g2_decap_8 FILLER_45_542 ();
 sg13g2_decap_8 FILLER_45_549 ();
 sg13g2_decap_8 FILLER_45_556 ();
 sg13g2_decap_8 FILLER_45_563 ();
 sg13g2_decap_8 FILLER_45_570 ();
 sg13g2_decap_8 FILLER_45_577 ();
 sg13g2_decap_8 FILLER_45_584 ();
 sg13g2_decap_8 FILLER_45_591 ();
 sg13g2_decap_8 FILLER_45_598 ();
 sg13g2_decap_8 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_612 ();
 sg13g2_decap_8 FILLER_45_619 ();
 sg13g2_decap_8 FILLER_45_626 ();
 sg13g2_decap_8 FILLER_45_633 ();
 sg13g2_decap_8 FILLER_45_640 ();
 sg13g2_decap_8 FILLER_45_647 ();
 sg13g2_decap_8 FILLER_45_654 ();
 sg13g2_decap_8 FILLER_45_661 ();
 sg13g2_decap_8 FILLER_45_668 ();
 sg13g2_decap_8 FILLER_45_675 ();
 sg13g2_decap_8 FILLER_45_682 ();
 sg13g2_decap_8 FILLER_45_689 ();
 sg13g2_decap_8 FILLER_45_696 ();
 sg13g2_decap_8 FILLER_45_703 ();
 sg13g2_decap_8 FILLER_45_710 ();
 sg13g2_decap_8 FILLER_45_717 ();
 sg13g2_decap_8 FILLER_45_724 ();
 sg13g2_decap_8 FILLER_45_731 ();
 sg13g2_decap_8 FILLER_45_738 ();
 sg13g2_decap_8 FILLER_45_745 ();
 sg13g2_decap_8 FILLER_45_752 ();
 sg13g2_decap_8 FILLER_45_759 ();
 sg13g2_decap_8 FILLER_45_766 ();
 sg13g2_decap_8 FILLER_45_773 ();
 sg13g2_decap_8 FILLER_45_780 ();
 sg13g2_decap_8 FILLER_45_787 ();
 sg13g2_decap_8 FILLER_45_794 ();
 sg13g2_decap_8 FILLER_45_801 ();
 sg13g2_decap_8 FILLER_45_808 ();
 sg13g2_decap_8 FILLER_45_815 ();
 sg13g2_decap_8 FILLER_45_822 ();
 sg13g2_decap_8 FILLER_45_829 ();
 sg13g2_decap_8 FILLER_45_836 ();
 sg13g2_decap_8 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_850 ();
 sg13g2_decap_8 FILLER_45_857 ();
 sg13g2_decap_8 FILLER_45_864 ();
 sg13g2_decap_8 FILLER_45_871 ();
 sg13g2_decap_8 FILLER_45_878 ();
 sg13g2_decap_8 FILLER_45_885 ();
 sg13g2_decap_8 FILLER_45_892 ();
 sg13g2_decap_8 FILLER_45_899 ();
 sg13g2_decap_8 FILLER_45_906 ();
 sg13g2_decap_8 FILLER_45_913 ();
 sg13g2_decap_8 FILLER_45_920 ();
 sg13g2_decap_8 FILLER_45_927 ();
 sg13g2_decap_8 FILLER_45_934 ();
 sg13g2_decap_8 FILLER_45_941 ();
 sg13g2_decap_8 FILLER_45_948 ();
 sg13g2_decap_8 FILLER_45_955 ();
 sg13g2_decap_8 FILLER_45_962 ();
 sg13g2_decap_8 FILLER_45_969 ();
 sg13g2_decap_8 FILLER_45_976 ();
 sg13g2_decap_8 FILLER_45_983 ();
 sg13g2_decap_8 FILLER_45_990 ();
 sg13g2_decap_8 FILLER_45_997 ();
 sg13g2_decap_8 FILLER_45_1004 ();
 sg13g2_decap_8 FILLER_45_1011 ();
 sg13g2_decap_8 FILLER_45_1018 ();
 sg13g2_decap_4 FILLER_45_1025 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_fill_1 FILLER_46_91 ();
 sg13g2_decap_4 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_180 ();
 sg13g2_fill_2 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_fill_2 FILLER_46_210 ();
 sg13g2_fill_1 FILLER_46_212 ();
 sg13g2_decap_8 FILLER_46_222 ();
 sg13g2_decap_8 FILLER_46_229 ();
 sg13g2_decap_4 FILLER_46_236 ();
 sg13g2_fill_2 FILLER_46_240 ();
 sg13g2_fill_2 FILLER_46_246 ();
 sg13g2_fill_1 FILLER_46_362 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_decap_8 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_decap_8 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_46_868 ();
 sg13g2_decap_8 FILLER_46_875 ();
 sg13g2_decap_8 FILLER_46_882 ();
 sg13g2_decap_8 FILLER_46_889 ();
 sg13g2_decap_8 FILLER_46_896 ();
 sg13g2_decap_8 FILLER_46_903 ();
 sg13g2_decap_8 FILLER_46_910 ();
 sg13g2_decap_8 FILLER_46_917 ();
 sg13g2_decap_8 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_46_931 ();
 sg13g2_decap_8 FILLER_46_938 ();
 sg13g2_decap_8 FILLER_46_945 ();
 sg13g2_decap_8 FILLER_46_952 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_decap_8 FILLER_46_966 ();
 sg13g2_decap_8 FILLER_46_973 ();
 sg13g2_decap_8 FILLER_46_980 ();
 sg13g2_decap_8 FILLER_46_987 ();
 sg13g2_decap_8 FILLER_46_994 ();
 sg13g2_decap_8 FILLER_46_1001 ();
 sg13g2_decap_8 FILLER_46_1008 ();
 sg13g2_decap_8 FILLER_46_1015 ();
 sg13g2_decap_8 FILLER_46_1022 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_4 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_95 ();
 sg13g2_decap_8 FILLER_47_101 ();
 sg13g2_decap_8 FILLER_47_108 ();
 sg13g2_decap_8 FILLER_47_115 ();
 sg13g2_fill_2 FILLER_47_122 ();
 sg13g2_decap_8 FILLER_47_142 ();
 sg13g2_decap_4 FILLER_47_149 ();
 sg13g2_fill_1 FILLER_47_153 ();
 sg13g2_decap_8 FILLER_47_167 ();
 sg13g2_decap_8 FILLER_47_174 ();
 sg13g2_decap_8 FILLER_47_181 ();
 sg13g2_decap_8 FILLER_47_188 ();
 sg13g2_decap_8 FILLER_47_195 ();
 sg13g2_decap_8 FILLER_47_202 ();
 sg13g2_decap_8 FILLER_47_209 ();
 sg13g2_decap_8 FILLER_47_216 ();
 sg13g2_decap_8 FILLER_47_223 ();
 sg13g2_decap_8 FILLER_47_230 ();
 sg13g2_decap_8 FILLER_47_237 ();
 sg13g2_decap_8 FILLER_47_244 ();
 sg13g2_fill_2 FILLER_47_251 ();
 sg13g2_fill_2 FILLER_47_257 ();
 sg13g2_fill_1 FILLER_47_259 ();
 sg13g2_decap_4 FILLER_47_270 ();
 sg13g2_fill_1 FILLER_47_274 ();
 sg13g2_fill_1 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_294 ();
 sg13g2_fill_2 FILLER_47_298 ();
 sg13g2_fill_1 FILLER_47_313 ();
 sg13g2_fill_1 FILLER_47_332 ();
 sg13g2_decap_8 FILLER_47_346 ();
 sg13g2_decap_8 FILLER_47_353 ();
 sg13g2_fill_2 FILLER_47_360 ();
 sg13g2_decap_8 FILLER_47_375 ();
 sg13g2_decap_8 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_47_389 ();
 sg13g2_fill_2 FILLER_47_396 ();
 sg13g2_fill_1 FILLER_47_398 ();
 sg13g2_fill_2 FILLER_47_412 ();
 sg13g2_decap_8 FILLER_47_423 ();
 sg13g2_decap_8 FILLER_47_430 ();
 sg13g2_decap_8 FILLER_47_437 ();
 sg13g2_decap_8 FILLER_47_444 ();
 sg13g2_decap_8 FILLER_47_451 ();
 sg13g2_decap_8 FILLER_47_458 ();
 sg13g2_decap_8 FILLER_47_465 ();
 sg13g2_decap_8 FILLER_47_472 ();
 sg13g2_decap_8 FILLER_47_479 ();
 sg13g2_decap_8 FILLER_47_486 ();
 sg13g2_decap_8 FILLER_47_493 ();
 sg13g2_decap_8 FILLER_47_500 ();
 sg13g2_decap_8 FILLER_47_507 ();
 sg13g2_decap_8 FILLER_47_514 ();
 sg13g2_decap_8 FILLER_47_521 ();
 sg13g2_decap_8 FILLER_47_528 ();
 sg13g2_decap_8 FILLER_47_535 ();
 sg13g2_decap_8 FILLER_47_542 ();
 sg13g2_decap_8 FILLER_47_549 ();
 sg13g2_decap_8 FILLER_47_556 ();
 sg13g2_decap_8 FILLER_47_563 ();
 sg13g2_decap_8 FILLER_47_570 ();
 sg13g2_decap_8 FILLER_47_577 ();
 sg13g2_decap_8 FILLER_47_584 ();
 sg13g2_decap_8 FILLER_47_591 ();
 sg13g2_decap_8 FILLER_47_598 ();
 sg13g2_decap_8 FILLER_47_605 ();
 sg13g2_decap_8 FILLER_47_612 ();
 sg13g2_decap_8 FILLER_47_619 ();
 sg13g2_decap_8 FILLER_47_626 ();
 sg13g2_decap_8 FILLER_47_633 ();
 sg13g2_decap_8 FILLER_47_640 ();
 sg13g2_decap_8 FILLER_47_647 ();
 sg13g2_decap_8 FILLER_47_654 ();
 sg13g2_decap_8 FILLER_47_661 ();
 sg13g2_decap_8 FILLER_47_668 ();
 sg13g2_decap_8 FILLER_47_675 ();
 sg13g2_decap_8 FILLER_47_682 ();
 sg13g2_decap_8 FILLER_47_689 ();
 sg13g2_decap_8 FILLER_47_696 ();
 sg13g2_decap_8 FILLER_47_703 ();
 sg13g2_decap_8 FILLER_47_710 ();
 sg13g2_decap_8 FILLER_47_717 ();
 sg13g2_decap_8 FILLER_47_724 ();
 sg13g2_decap_8 FILLER_47_731 ();
 sg13g2_decap_8 FILLER_47_738 ();
 sg13g2_decap_8 FILLER_47_745 ();
 sg13g2_decap_8 FILLER_47_752 ();
 sg13g2_decap_8 FILLER_47_759 ();
 sg13g2_decap_8 FILLER_47_766 ();
 sg13g2_decap_8 FILLER_47_773 ();
 sg13g2_decap_8 FILLER_47_780 ();
 sg13g2_decap_8 FILLER_47_787 ();
 sg13g2_decap_8 FILLER_47_794 ();
 sg13g2_decap_8 FILLER_47_801 ();
 sg13g2_decap_8 FILLER_47_808 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_decap_8 FILLER_47_843 ();
 sg13g2_decap_8 FILLER_47_850 ();
 sg13g2_decap_8 FILLER_47_857 ();
 sg13g2_decap_8 FILLER_47_864 ();
 sg13g2_decap_8 FILLER_47_871 ();
 sg13g2_decap_8 FILLER_47_878 ();
 sg13g2_decap_8 FILLER_47_885 ();
 sg13g2_decap_8 FILLER_47_892 ();
 sg13g2_decap_8 FILLER_47_899 ();
 sg13g2_decap_8 FILLER_47_906 ();
 sg13g2_decap_8 FILLER_47_913 ();
 sg13g2_decap_8 FILLER_47_920 ();
 sg13g2_decap_8 FILLER_47_927 ();
 sg13g2_decap_8 FILLER_47_934 ();
 sg13g2_decap_8 FILLER_47_941 ();
 sg13g2_decap_8 FILLER_47_948 ();
 sg13g2_decap_8 FILLER_47_955 ();
 sg13g2_decap_8 FILLER_47_962 ();
 sg13g2_decap_8 FILLER_47_969 ();
 sg13g2_decap_8 FILLER_47_976 ();
 sg13g2_decap_8 FILLER_47_983 ();
 sg13g2_decap_8 FILLER_47_990 ();
 sg13g2_decap_8 FILLER_47_997 ();
 sg13g2_decap_8 FILLER_47_1004 ();
 sg13g2_decap_8 FILLER_47_1011 ();
 sg13g2_decap_8 FILLER_47_1018 ();
 sg13g2_decap_4 FILLER_47_1025 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_4 FILLER_48_318 ();
 sg13g2_fill_2 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_333 ();
 sg13g2_decap_8 FILLER_48_340 ();
 sg13g2_decap_8 FILLER_48_347 ();
 sg13g2_decap_8 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_361 ();
 sg13g2_decap_8 FILLER_48_368 ();
 sg13g2_decap_8 FILLER_48_375 ();
 sg13g2_decap_8 FILLER_48_382 ();
 sg13g2_decap_8 FILLER_48_389 ();
 sg13g2_decap_8 FILLER_48_396 ();
 sg13g2_decap_8 FILLER_48_403 ();
 sg13g2_decap_8 FILLER_48_410 ();
 sg13g2_decap_8 FILLER_48_417 ();
 sg13g2_decap_8 FILLER_48_424 ();
 sg13g2_decap_8 FILLER_48_431 ();
 sg13g2_decap_8 FILLER_48_438 ();
 sg13g2_decap_8 FILLER_48_445 ();
 sg13g2_decap_8 FILLER_48_452 ();
 sg13g2_decap_8 FILLER_48_459 ();
 sg13g2_decap_8 FILLER_48_466 ();
 sg13g2_decap_8 FILLER_48_473 ();
 sg13g2_decap_8 FILLER_48_480 ();
 sg13g2_decap_8 FILLER_48_487 ();
 sg13g2_decap_8 FILLER_48_494 ();
 sg13g2_decap_8 FILLER_48_501 ();
 sg13g2_decap_8 FILLER_48_508 ();
 sg13g2_decap_8 FILLER_48_515 ();
 sg13g2_decap_8 FILLER_48_522 ();
 sg13g2_decap_8 FILLER_48_529 ();
 sg13g2_decap_8 FILLER_48_536 ();
 sg13g2_decap_8 FILLER_48_543 ();
 sg13g2_decap_8 FILLER_48_550 ();
 sg13g2_decap_8 FILLER_48_557 ();
 sg13g2_decap_8 FILLER_48_564 ();
 sg13g2_decap_8 FILLER_48_571 ();
 sg13g2_decap_8 FILLER_48_578 ();
 sg13g2_decap_8 FILLER_48_585 ();
 sg13g2_decap_8 FILLER_48_592 ();
 sg13g2_decap_8 FILLER_48_599 ();
 sg13g2_decap_8 FILLER_48_606 ();
 sg13g2_decap_8 FILLER_48_613 ();
 sg13g2_decap_8 FILLER_48_620 ();
 sg13g2_decap_8 FILLER_48_627 ();
 sg13g2_decap_8 FILLER_48_634 ();
 sg13g2_decap_8 FILLER_48_641 ();
 sg13g2_decap_8 FILLER_48_648 ();
 sg13g2_decap_8 FILLER_48_655 ();
 sg13g2_decap_8 FILLER_48_662 ();
 sg13g2_decap_8 FILLER_48_669 ();
 sg13g2_decap_8 FILLER_48_676 ();
 sg13g2_decap_8 FILLER_48_683 ();
 sg13g2_decap_8 FILLER_48_690 ();
 sg13g2_decap_8 FILLER_48_697 ();
 sg13g2_decap_8 FILLER_48_704 ();
 sg13g2_decap_8 FILLER_48_711 ();
 sg13g2_decap_8 FILLER_48_718 ();
 sg13g2_decap_8 FILLER_48_725 ();
 sg13g2_decap_8 FILLER_48_732 ();
 sg13g2_decap_8 FILLER_48_739 ();
 sg13g2_decap_8 FILLER_48_746 ();
 sg13g2_decap_8 FILLER_48_753 ();
 sg13g2_decap_8 FILLER_48_760 ();
 sg13g2_decap_8 FILLER_48_767 ();
 sg13g2_decap_8 FILLER_48_774 ();
 sg13g2_decap_8 FILLER_48_781 ();
 sg13g2_decap_8 FILLER_48_788 ();
 sg13g2_decap_8 FILLER_48_795 ();
 sg13g2_decap_8 FILLER_48_802 ();
 sg13g2_decap_8 FILLER_48_809 ();
 sg13g2_decap_8 FILLER_48_816 ();
 sg13g2_decap_8 FILLER_48_823 ();
 sg13g2_decap_8 FILLER_48_830 ();
 sg13g2_decap_8 FILLER_48_837 ();
 sg13g2_decap_8 FILLER_48_844 ();
 sg13g2_decap_8 FILLER_48_851 ();
 sg13g2_decap_8 FILLER_48_858 ();
 sg13g2_decap_8 FILLER_48_865 ();
 sg13g2_decap_8 FILLER_48_872 ();
 sg13g2_decap_8 FILLER_48_879 ();
 sg13g2_decap_8 FILLER_48_886 ();
 sg13g2_decap_8 FILLER_48_893 ();
 sg13g2_decap_8 FILLER_48_900 ();
 sg13g2_decap_8 FILLER_48_907 ();
 sg13g2_decap_8 FILLER_48_914 ();
 sg13g2_decap_8 FILLER_48_921 ();
 sg13g2_decap_8 FILLER_48_928 ();
 sg13g2_decap_8 FILLER_48_935 ();
 sg13g2_decap_8 FILLER_48_942 ();
 sg13g2_decap_8 FILLER_48_949 ();
 sg13g2_decap_8 FILLER_48_956 ();
 sg13g2_decap_8 FILLER_48_963 ();
 sg13g2_decap_8 FILLER_48_970 ();
 sg13g2_decap_8 FILLER_48_977 ();
 sg13g2_decap_8 FILLER_48_984 ();
 sg13g2_decap_8 FILLER_48_991 ();
 sg13g2_decap_8 FILLER_48_998 ();
 sg13g2_decap_8 FILLER_48_1005 ();
 sg13g2_decap_8 FILLER_48_1012 ();
 sg13g2_decap_8 FILLER_48_1019 ();
 sg13g2_fill_2 FILLER_48_1026 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_8 FILLER_49_497 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_882 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_decap_8 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_973 ();
 sg13g2_decap_8 FILLER_49_980 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
 assign uo_out[1] = net19;
 assign uo_out[2] = net20;
 assign uo_out[3] = net21;
 assign uo_out[4] = net22;
 assign uo_out[5] = net23;
 assign uo_out[6] = net24;
 assign uo_out[7] = net25;
endmodule
